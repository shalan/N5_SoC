* NGSPICE file created from apb_sys_0.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt apb_sys_0 HADDR[0] HADDR[10] HADDR[11] HADDR[12] HADDR[13] HADDR[14] HADDR[15]
+ HADDR[16] HADDR[17] HADDR[18] HADDR[19] HADDR[1] HADDR[20] HADDR[21] HADDR[22] HADDR[23]
+ HADDR[24] HADDR[25] HADDR[26] HADDR[27] HADDR[28] HADDR[29] HADDR[2] HADDR[30] HADDR[31]
+ HADDR[3] HADDR[4] HADDR[5] HADDR[6] HADDR[7] HADDR[8] HADDR[9] HCLK HRDATA[0] HRDATA[10]
+ HRDATA[11] HRDATA[12] HRDATA[13] HRDATA[14] HRDATA[15] HRDATA[16] HRDATA[17] HRDATA[18]
+ HRDATA[19] HRDATA[1] HRDATA[20] HRDATA[21] HRDATA[22] HRDATA[23] HRDATA[24] HRDATA[25]
+ HRDATA[26] HRDATA[27] HRDATA[28] HRDATA[29] HRDATA[2] HRDATA[30] HRDATA[31] HRDATA[3]
+ HRDATA[4] HRDATA[5] HRDATA[6] HRDATA[7] HRDATA[8] HRDATA[9] HREADY HREADYOUT HRESETn
+ HSEL HTRANS[0] HTRANS[1] HWDATA[0] HWDATA[10] HWDATA[11] HWDATA[12] HWDATA[13] HWDATA[14]
+ HWDATA[15] HWDATA[16] HWDATA[17] HWDATA[18] HWDATA[19] HWDATA[1] HWDATA[20] HWDATA[21]
+ HWDATA[22] HWDATA[23] HWDATA[24] HWDATA[25] HWDATA[26] HWDATA[27] HWDATA[28] HWDATA[29]
+ HWDATA[2] HWDATA[30] HWDATA[31] HWDATA[3] HWDATA[4] HWDATA[5] HWDATA[6] HWDATA[7]
+ HWDATA[8] HWDATA[9] HWRITE IRQ[0] IRQ[10] IRQ[11] IRQ[12] IRQ[13] IRQ[14] IRQ[15]
+ IRQ[1] IRQ[2] IRQ[3] IRQ[4] IRQ[5] IRQ[6] IRQ[7] IRQ[8] IRQ[9] MSI_S2 MSI_S3 MSO_S2
+ MSO_S3 RsRx_S0 RsRx_S1 RsTx_S0 RsTx_S1 SCLK_S2 SCLK_S3 SSn_S2 SSn_S3 pwm_S6 pwm_S7
+ scl_i_S4 scl_i_S5 scl_o_S4 scl_o_S5 scl_oen_o_S4 scl_oen_o_S5 sda_i_S4 sda_i_S5
+ sda_o_S4 sda_o_S5 sda_oen_o_S4 sda_oen_o_S5 VPWR VGND
XANTENNA__18243__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18869_ _18868_/Y VGND VGND VPWR VPWR _18869_/X sky130_fd_sc_hd__buf_2
X_20900_ _20900_/A _20900_/B VGND VGND VPWR VPWR _20901_/A sky130_fd_sc_hd__or2_4
XANTENNA__13615__A _14645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21880_ _21245_/A VGND VGND VPWR VPWR _21886_/A sky130_fd_sc_hd__buf_2
XFILLER_55_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20831_ _20830_/X VGND VGND VPWR VPWR _24032_/D sky130_fd_sc_hd__inv_2
XFILLER_36_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24992__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22647__B _22644_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20762_ _20761_/X VGND VGND VPWR VPWR _20767_/B sky130_fd_sc_hd__inv_2
XANTENNA__24921__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23550_ _23550_/CLK _19946_/X VGND VGND VPWR VPWR _19945_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_35_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22501_ _12023_/Y _13533_/B _12092_/Y _12060_/B VGND VGND VPWR VPWR _22501_/X sky130_fd_sc_hd__o22a_4
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24239__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23481_ _23496_/CLK _20136_/X VGND VGND VPWR VPWR _23481_/Q sky130_fd_sc_hd__dfxtp_4
X_20693_ _20692_/X VGND VGND VPWR VPWR _24000_/D sky130_fd_sc_hd__inv_2
XFILLER_50_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_13_0_HCLK_A clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22432_ _22714_/A _22430_/X _21438_/X _22431_/X VGND VGND VPWR VPWR _22433_/A sky130_fd_sc_hd__o22a_4
XFILLER_17_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25220_ _25043_/CLK _25220_/D HRESETn VGND VGND VPWR VPWR _25220_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16309__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22645__A3 _22130_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22363_ _22070_/X _22363_/B VGND VGND VPWR VPWR _22363_/X sky130_fd_sc_hd__or2_4
XANTENNA__21853__A1 _24707_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12594__B2 _24846_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25151_ _24109_/CLK _14347_/X HRESETn VGND VGND VPWR VPWR _25151_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21314_ _21314_/A _21314_/B VGND VGND VPWR VPWR _21314_/X sky130_fd_sc_hd__or2_4
X_24102_ _24102_/CLK _12154_/X HRESETn VGND VGND VPWR VPWR _12152_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21279__A _21859_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25082_ _24376_/CLK _14585_/X HRESETn VGND VGND VPWR VPWR _14558_/A sky130_fd_sc_hd__dfrtp_4
X_22294_ _22294_/A _22927_/A VGND VGND VPWR VPWR _22297_/B sky130_fd_sc_hd__or2_4
XFILLER_50_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17476__B _17449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24033_ _24033_/CLK _20835_/Y HRESETn VGND VGND VPWR VPWR _13656_/A sky130_fd_sc_hd__dfrtp_4
X_21245_ _21245_/A _20165_/Y VGND VGND VPWR VPWR _21245_/X sky130_fd_sc_hd__or2_4
XANTENNA__25098__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21176_ _21184_/A _21176_/B VGND VGND VPWR VPWR _21176_/X sky130_fd_sc_hd__or2_4
XFILLER_132_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25027__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20127_ _20127_/A VGND VGND VPWR VPWR _20140_/A sky130_fd_sc_hd__inv_2
XFILLER_137_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18234__B1 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20058_ _20056_/Y _20057_/X _19794_/X _20057_/X VGND VGND VPWR VPWR _23511_/D sky130_fd_sc_hd__a2bb2o_4
X_24935_ _24248_/CLK _15493_/X HRESETn VGND VGND VPWR VPWR _12052_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14415__A1_N _14128_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11900_ _11900_/A _11871_/Y VGND VGND VPWR VPWR _11901_/A sky130_fd_sc_hd__and2_4
XANTENNA__22581__A2 _22578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12880_ _12880_/A _12880_/B VGND VGND VPWR VPWR _12881_/C sky130_fd_sc_hd__or2_4
XFILLER_73_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24866_ _24847_/CLK _15727_/X HRESETn VGND VGND VPWR VPWR _12539_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_22_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22838__A _23021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_128_0_HCLK clkbuf_7_64_0_HCLK/X VGND VGND VPWR VPWR _23718_/CLK sky130_fd_sc_hd__clkbuf_1
X_11831_ _11831_/A VGND VGND VPWR VPWR _11831_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23817_ _23832_/CLK _23817_/D VGND VGND VPWR VPWR _23817_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _24832_/CLK _15875_/X HRESETn VGND VGND VPWR VPWR _24797_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16836__A _24412_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15740__A _15740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14550_ _25086_/Q _14066_/X _14060_/X VGND VGND VPWR VPWR _25086_/D sky130_fd_sc_hd__a21bo_4
XFILLER_54_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19212__A _16442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24662__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11759_/Y _11760_/X _11761_/X _11760_/X VGND VGND VPWR VPWR _11762_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16548__B1 _16285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ _23828_/CLK _23748_/D VGND VGND VPWR VPWR _17946_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13497_/Y VGND VGND VPWR VPWR _13501_/X sky130_fd_sc_hd__buf_2
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14481_/A VGND VGND VPWR VPWR _14481_/X sky130_fd_sc_hd__buf_2
X_11693_ _25270_/Q VGND VGND VPWR VPWR _13729_/A sky130_fd_sc_hd__inv_2
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23679_ _23398_/CLK _19575_/X VGND VGND VPWR VPWR _23679_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15220__B1 _15174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16219_/Y _16217_/X _15962_/X _16217_/X VGND VGND VPWR VPWR _16220_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _13196_/Y _13431_/X _25314_/Q _13195_/X VGND VGND VPWR VPWR _25314_/D sky130_fd_sc_hd__o22a_4
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25418_ _25411_/CLK _12632_/Y HRESETn VGND VGND VPWR VPWR _12592_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16151_ _22183_/A VGND VGND VPWR VPWR _16151_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12585__B2 _12584_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13363_ _13395_/A _13363_/B VGND VGND VPWR VPWR _13363_/X sky130_fd_sc_hd__or2_4
XANTENNA__21844__B2 _17416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25349_ _23370_/CLK _13024_/X HRESETn VGND VGND VPWR VPWR _25349_/Q sky130_fd_sc_hd__dfrtp_4
X_15102_ _24591_/Q VGND VGND VPWR VPWR _15102_/Y sky130_fd_sc_hd__inv_2
X_12314_ _12314_/A VGND VGND VPWR VPWR _12988_/A sky130_fd_sc_hd__inv_2
X_16082_ _11739_/A _15668_/X _15927_/X _24700_/Q _16081_/X VGND VGND VPWR VPWR _24700_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13294_ _13366_/A _13285_/X _13293_/X VGND VGND VPWR VPWR _13294_/X sky130_fd_sc_hd__and3_4
XFILLER_114_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15033_ _15024_/X _15033_/B _15029_/X _15032_/X VGND VGND VPWR VPWR _15055_/A sky130_fd_sc_hd__or4_4
X_19910_ _19909_/X VGND VGND VPWR VPWR _19923_/A sky130_fd_sc_hd__inv_2
XANTENNA__15187__A _15187_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12245_ _12244_/Y _24758_/Q _12244_/Y _24758_/Q VGND VGND VPWR VPWR _12245_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12604__A _12604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25450__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12176_ _14329_/A _12173_/Y _11867_/X _12173_/Y VGND VGND VPWR VPWR _12176_/X sky130_fd_sc_hd__a2bb2o_4
X_19841_ _19841_/A VGND VGND VPWR VPWR _19841_/X sky130_fd_sc_hd__buf_2
XFILLER_123_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15915__A _25289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16984_ _24712_/Q _16983_/A _16051_/Y _17038_/A VGND VGND VPWR VPWR _16989_/B sky130_fd_sc_hd__o22a_4
X_19772_ _19770_/Y _19766_/X _19771_/X _19751_/Y VGND VGND VPWR VPWR _19772_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12250__A1_N _12249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15935_ _15894_/A VGND VGND VPWR VPWR _15935_/X sky130_fd_sc_hd__buf_2
X_18723_ _18694_/X _18703_/X _18672_/Y VGND VGND VPWR VPWR _18724_/C sky130_fd_sc_hd__o21a_4
Xclkbuf_7_24_0_HCLK clkbuf_7_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_49_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13435__A _13233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22572__A2 _22525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18654_ _24141_/Q VGND VGND VPWR VPWR _18654_/Y sky130_fd_sc_hd__inv_2
X_15866_ _15850_/X _15857_/X _15714_/X _24802_/Q _15864_/X VGND VGND VPWR VPWR _24802_/D
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_7_87_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_87_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14817_ _25039_/Q _14816_/X _14817_/C VGND VGND VPWR VPWR _14817_/X sky130_fd_sc_hd__or3_4
X_17605_ _17605_/A _17604_/Y VGND VGND VPWR VPWR _17607_/B sky130_fd_sc_hd__or2_4
XFILLER_40_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18585_ _18475_/C _18592_/A VGND VGND VPWR VPWR _18585_/X sky130_fd_sc_hd__or2_4
X_15797_ _15817_/A VGND VGND VPWR VPWR _15829_/A sky130_fd_sc_hd__inv_2
XFILLER_17_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12265__A1_N _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17536_ _11798_/Y _17565_/A _11798_/Y _17565_/A VGND VGND VPWR VPWR _17536_/X sky130_fd_sc_hd__a2bb2o_4
X_14748_ _14676_/A VGND VGND VPWR VPWR _14749_/A sky130_fd_sc_hd__buf_2
XFILLER_127_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16566__A1_N _16565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23987__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17200__B2 _17199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24332__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17467_ _24194_/Q VGND VGND VPWR VPWR _17467_/Y sky130_fd_sc_hd__inv_2
X_14679_ _14679_/A VGND VGND VPWR VPWR _21371_/A sky130_fd_sc_hd__buf_2
XANTENNA__18961__A _16442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16418_ _24581_/Q VGND VGND VPWR VPWR _16418_/Y sky130_fd_sc_hd__inv_2
X_19206_ _16781_/X VGND VGND VPWR VPWR _19206_/X sky130_fd_sc_hd__buf_2
X_17398_ _23980_/Q _17398_/B VGND VGND VPWR VPWR _17399_/B sky130_fd_sc_hd__or2_4
XANTENNA__22483__A _22186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19137_ _19130_/A VGND VGND VPWR VPWR _19137_/X sky130_fd_sc_hd__buf_2
XFILLER_125_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21835__A1 _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16349_ _22273_/A VGND VGND VPWR VPWR _16349_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25538__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19068_ _19062_/Y VGND VGND VPWR VPWR _19068_/X sky130_fd_sc_hd__buf_2
XANTENNA__23037__B1 _24865_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18019_ _18019_/A VGND VGND VPWR VPWR _18019_/X sky130_fd_sc_hd__buf_2
XFILLER_114_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12514__A _12514_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21030_ _21030_/A VGND VGND VPWR VPWR _21030_/X sky130_fd_sc_hd__buf_2
XANTENNA__25191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21827__A _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15760__A1_N _12536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16519__A1_N _16518_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11839__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22981_ _12285_/C _22980_/X _16900_/A _22906_/X VGND VGND VPWR VPWR _22981_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12500__A1 _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24720_ _24720_/CLK _16032_/X HRESETn VGND VGND VPWR VPWR _24720_/Q sky130_fd_sc_hd__dfrtp_4
X_21932_ _21927_/X _21931_/X _18298_/X VGND VGND VPWR VPWR _21932_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21562__A _16453_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24651_ _24162_/CLK _24651_/D HRESETn VGND VGND VPWR VPWR _22809_/A sky130_fd_sc_hd__dfrtp_4
X_21863_ _23034_/A VGND VGND VPWR VPWR _21863_/X sky130_fd_sc_hd__buf_2
XFILLER_103_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19716__B1 _19715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23602_ _23618_/CLK _19809_/X VGND VGND VPWR VPWR _19807_/A sky130_fd_sc_hd__dfxtp_4
X_20814_ _20863_/A VGND VGND VPWR VPWR _20814_/X sky130_fd_sc_hd__buf_2
X_21794_ _21460_/A _21792_/X _21794_/C VGND VGND VPWR VPWR _21794_/X sky130_fd_sc_hd__and3_4
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24582_ _24572_/CLK _16417_/X HRESETn VGND VGND VPWR VPWR _24582_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24073__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23533_ _23533_/CLK _23533_/D VGND VGND VPWR VPWR _23533_/Q sky130_fd_sc_hd__dfxtp_4
X_20745_ _20772_/C VGND VGND VPWR VPWR _20745_/Y sky130_fd_sc_hd__inv_2
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24002__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20676_ _20724_/A VGND VGND VPWR VPWR _20676_/X sky130_fd_sc_hd__buf_2
XANTENNA__15753__A1 _15749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23276__B1 _24733_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23464_ _23496_/CLK _23464_/D VGND VGND VPWR VPWR _20179_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22393__A _22523_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25203_ _25199_/CLK _25203_/D HRESETn VGND VGND VPWR VPWR _14100_/A sky130_fd_sc_hd__dfrtp_4
X_22415_ _25362_/Q _22288_/X _22414_/X VGND VGND VPWR VPWR _22415_/X sky130_fd_sc_hd__a21o_4
X_23395_ _23580_/CLK _23395_/D VGND VGND VPWR VPWR _20358_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__25279__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25134_ _23959_/CLK _14401_/X HRESETn VGND VGND VPWR VPWR _14399_/A sky130_fd_sc_hd__dfrtp_4
X_22346_ _21455_/A _22346_/B VGND VGND VPWR VPWR _22346_/X sky130_fd_sc_hd__or2_4
XANTENNA__13516__B1 _13515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12319__B2 _12318_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22277_ _22962_/A VGND VGND VPWR VPWR _23281_/A sky130_fd_sc_hd__buf_2
XFILLER_124_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25065_ _23826_/CLK _14642_/X HRESETn VGND VGND VPWR VPWR _13630_/A sky130_fd_sc_hd__dfrtp_4
X_12030_ _11989_/Y _12029_/X _25481_/Q _12029_/X VGND VGND VPWR VPWR _12030_/X sky130_fd_sc_hd__a2bb2o_4
X_21228_ _21377_/A VGND VGND VPWR VPWR _21250_/A sky130_fd_sc_hd__buf_2
X_24016_ _24018_/CLK _20765_/Y HRESETn VGND VGND VPWR VPWR _13119_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_105_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21159_ _21148_/X _21159_/B _21158_/X VGND VGND VPWR VPWR _21208_/C sky130_fd_sc_hd__and3_4
XFILLER_104_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18655__A1_N _16613_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13981_ _14002_/A VGND VGND VPWR VPWR _13982_/A sky130_fd_sc_hd__buf_2
XFILLER_111_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15720_ _12582_/Y _15718_/X _11754_/X _15718_/X VGND VGND VPWR VPWR _24870_/D sky130_fd_sc_hd__a2bb2o_4
X_12932_ _12799_/X _12931_/X VGND VGND VPWR VPWR _12933_/A sky130_fd_sc_hd__or2_4
XFILLER_24_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24918_ _25433_/CLK _24918_/D HRESETn VGND VGND VPWR VPWR _11726_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__24843__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15651_ _15643_/Y _15646_/X _15647_/X _21008_/B _15650_/X VGND VGND VPWR VPWR _24879_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_2_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12863_ _12855_/X _12862_/X VGND VGND VPWR VPWR _12863_/X sky130_fd_sc_hd__or2_4
X_24849_ _23370_/CLK _24849_/D HRESETn VGND VGND VPWR VPWR _12542_/A sky130_fd_sc_hd__dfrtp_4
X_14602_ _13769_/Y VGND VGND VPWR VPWR _14602_/X sky130_fd_sc_hd__buf_2
XANTENNA__22287__B _22286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11814_ _11811_/Y _11805_/X _11813_/X _11805_/X VGND VGND VPWR VPWR _11814_/X sky130_fd_sc_hd__a2bb2o_4
X_18370_ _18370_/A _18370_/B _14339_/A _12157_/X VGND VGND VPWR VPWR _18371_/A sky130_fd_sc_hd__or4_4
X_15582_ _15579_/Y _15575_/X _11771_/X _15581_/X VGND VGND VPWR VPWR _15582_/X sky130_fd_sc_hd__a2bb2o_4
X_12794_ _12810_/A _12792_/Y _12959_/A _24777_/Q VGND VGND VPWR VPWR _12804_/A sky130_fd_sc_hd__a2bb2o_4
XPHY_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17203_/Y _17321_/B VGND VGND VPWR VPWR _17321_/X sky130_fd_sc_hd__or2_4
XFILLER_42_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14533_ _23951_/Q _14532_/X _25101_/Q _14517_/A VGND VGND VPWR VPWR _14533_/X sky130_fd_sc_hd__o22a_4
XFILLER_42_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _25537_/Q VGND VGND VPWR VPWR _11745_/Y sky130_fd_sc_hd__inv_2
XPHY_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17252_/A _17252_/B _17252_/C _17220_/Y VGND VGND VPWR VPWR _17252_/X sky130_fd_sc_hd__or4_4
X_14464_ _14463_/Y _14459_/X _14403_/X _14459_/X VGND VGND VPWR VPWR _25112_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _25273_/Q VGND VGND VPWR VPWR _13685_/A sky130_fd_sc_hd__inv_2
XFILLER_30_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ _16202_/Y _16200_/X _11764_/X _16200_/X VGND VGND VPWR VPWR _24659_/D sky130_fd_sc_hd__a2bb2o_4
X_13415_ _13297_/X _13407_/X _13415_/C VGND VGND VPWR VPWR _13415_/X sky130_fd_sc_hd__and3_4
XFILLER_127_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21817__A1 _20329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17183_ _22860_/A _24346_/Q _16318_/Y _17254_/A VGND VGND VPWR VPWR _17183_/X sky130_fd_sc_hd__o22a_4
XFILLER_122_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14395_ _15986_/A VGND VGND VPWR VPWR _14395_/X sky130_fd_sc_hd__buf_2
X_16134_ _16133_/Y _16131_/X _11809_/X _16131_/X VGND VGND VPWR VPWR _24681_/D sky130_fd_sc_hd__a2bb2o_4
X_13346_ _13309_/A _13344_/X _13345_/X VGND VGND VPWR VPWR _13350_/B sky130_fd_sc_hd__and3_4
XANTENNA__22490__B2 _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16065_ _16063_/Y _16060_/X _16064_/X _16060_/X VGND VGND VPWR VPWR _16065_/X sky130_fd_sc_hd__a2bb2o_4
X_13277_ _13225_/A VGND VGND VPWR VPWR _13316_/A sky130_fd_sc_hd__buf_2
XANTENNA__12334__A _24809_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15016_ _25022_/Q _15015_/Y _15283_/A _24434_/Q VGND VGND VPWR VPWR _15016_/X sky130_fd_sc_hd__a2bb2o_4
X_12228_ _24752_/Q VGND VGND VPWR VPWR _12228_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18446__B1 _16189_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20752__A1_N _20743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19824_ _19836_/A VGND VGND VPWR VPWR _19824_/X sky130_fd_sc_hd__buf_2
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19117__A _16786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15645__A _15648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12159_ _20965_/B VGND VGND VPWR VPWR _12159_/X sky130_fd_sc_hd__buf_2
XFILLER_81_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19755_ HWDATA[6] VGND VGND VPWR VPWR _19755_/X sky130_fd_sc_hd__buf_2
X_16967_ _16967_/A VGND VGND VPWR VPWR _17035_/A sky130_fd_sc_hd__inv_2
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18706_ _18669_/A VGND VGND VPWR VPWR _18733_/A sky130_fd_sc_hd__inv_2
X_15918_ _13588_/X _15693_/Y _15915_/X _15917_/Y VGND VGND VPWR VPWR _15918_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24584__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16898_ _16898_/A VGND VGND VPWR VPWR _16898_/X sky130_fd_sc_hd__buf_2
X_19686_ _19682_/Y _19685_/X _19664_/X _19685_/X VGND VGND VPWR VPWR _19686_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15849_ _15669_/X _15713_/A _15845_/X _12980_/A _15848_/X VGND VGND VPWR VPWR _24804_/D
+ sky130_fd_sc_hd__a32o_4
X_18637_ _24130_/Q VGND VGND VPWR VPWR _18757_/A sky130_fd_sc_hd__inv_2
XANTENNA__24513__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_111_0_HCLK clkbuf_7_55_0_HCLK/X VGND VGND VPWR VPWR _24035_/CLK sky130_fd_sc_hd__clkbuf_1
X_18568_ _18471_/Y _18566_/X _18567_/Y VGND VGND VPWR VPWR _18568_/X sky130_fd_sc_hd__o21a_4
XFILLER_91_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_174_0_HCLK clkbuf_7_87_0_HCLK/X VGND VGND VPWR VPWR _24930_/CLK sky130_fd_sc_hd__clkbuf_1
X_17519_ _24280_/Q VGND VGND VPWR VPWR _17662_/B sky130_fd_sc_hd__inv_2
XFILLER_36_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18499_ _18456_/A _18497_/X _18498_/X _18493_/B VGND VGND VPWR VPWR _18500_/A sky130_fd_sc_hd__a211o_4
XFILLER_127_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20530_ _17420_/A _20530_/B VGND VGND VPWR VPWR _23955_/D sky130_fd_sc_hd__and2_4
XFILLER_138_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23258__B1 _22090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20461_ _24063_/D VGND VGND VPWR VPWR _20461_/X sky130_fd_sc_hd__buf_2
XANTENNA__23102__A _21418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22200_ _22200_/A _19849_/Y VGND VGND VPWR VPWR _22202_/B sky130_fd_sc_hd__or2_4
XANTENNA__25372__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22481__A1 _22476_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23180_ _23143_/A _23180_/B VGND VGND VPWR VPWR _23190_/B sky130_fd_sc_hd__and2_4
X_20392_ _20383_/X _20379_/X _11862_/A _23381_/Q _20381_/X VGND VGND VPWR VPWR _20392_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22481__B2 _22480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22131_ _23306_/A _22122_/X _22127_/X _22130_/X VGND VGND VPWR VPWR _22132_/B sky130_fd_sc_hd__a211o_4
XANTENNA__25301__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23025__A3 _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22062_ _14682_/B _22062_/B VGND VGND VPWR VPWR _22062_/X sky130_fd_sc_hd__or2_4
XFILLER_47_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21013_ _12095_/A VGND VGND VPWR VPWR _21014_/A sky130_fd_sc_hd__buf_2
XANTENNA__15555__A _21154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22536__A2 _22534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22964_ _22964_/A _23140_/B VGND VGND VPWR VPWR _22964_/X sky130_fd_sc_hd__or2_4
XFILLER_83_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21292__A _21071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24703_ _24318_/CLK _16076_/X HRESETn VGND VGND VPWR VPWR _16075_/A sky130_fd_sc_hd__dfrtp_4
X_21915_ _21942_/A _21915_/B VGND VGND VPWR VPWR _21915_/X sky130_fd_sc_hd__or2_4
XANTENNA__24254__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_70_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_70_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16386__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22895_ _22895_/A _22472_/B VGND VGND VPWR VPWR _22895_/X sky130_fd_sc_hd__or2_4
XANTENNA__13803__A _15986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24634_ _24654_/CLK _16269_/X HRESETn VGND VGND VPWR VPWR _16268_/A sky130_fd_sc_hd__dfrtp_4
X_21846_ _12113_/Y _13496_/B _18379_/Y _12072_/D VGND VGND VPWR VPWR _21846_/X sky130_fd_sc_hd__o22a_4
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24565_ _24557_/CLK _16462_/X HRESETn VGND VGND VPWR VPWR _24565_/Q sky130_fd_sc_hd__dfrtp_4
X_21777_ _21759_/X _21776_/X _21821_/A VGND VGND VPWR VPWR _21777_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12419__A _12277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23516_ _23516_/CLK _20046_/X VGND VGND VPWR VPWR _20042_/A sky130_fd_sc_hd__dfxtp_4
X_20728_ _20728_/A VGND VGND VPWR VPWR _20728_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15726__A1 _15548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24496_ _24496_/CLK _24496_/D HRESETn VGND VGND VPWR VPWR _24496_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23447_ _23798_/CLK _23447_/D VGND VGND VPWR VPWR _20223_/A sky130_fd_sc_hd__dfxtp_4
X_20659_ _14226_/Y _20604_/Y _20619_/A _20658_/Y VGND VGND VPWR VPWR _20659_/X sky130_fd_sc_hd__a211o_4
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18106__A _18217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13200_ _13199_/Y VGND VGND VPWR VPWR _13200_/X sky130_fd_sc_hd__buf_2
XANTENNA__17479__A1 _21504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14180_ _14179_/X VGND VGND VPWR VPWR _25198_/D sky130_fd_sc_hd__inv_2
X_23378_ _23377_/CLK _20401_/X VGND VGND VPWR VPWR _23378_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25042__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13131_ _20728_/A _13131_/B VGND VGND VPWR VPWR _13132_/B sky130_fd_sc_hd__or2_4
XFILLER_137_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25117_ _25101_/CLK _14451_/X HRESETn VGND VGND VPWR VPWR _14182_/A sky130_fd_sc_hd__dfstp_4
X_22329_ _21942_/A _22329_/B VGND VGND VPWR VPWR _22329_/X sky130_fd_sc_hd__or2_4
XFILLER_136_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22224__A1 _21260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18428__B1 _22089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13062_ _13049_/A _13062_/B _13062_/C VGND VGND VPWR VPWR _13062_/X sky130_fd_sc_hd__and3_4
XANTENNA__21467__A _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25048_ _23494_/CLK _14759_/Y HRESETn VGND VGND VPWR VPWR _14679_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12013_ _11990_/Y _11997_/B _11997_/Y _12012_/X VGND VGND VPWR VPWR _12013_/X sky130_fd_sc_hd__a211o_4
X_17870_ _17867_/A _17867_/B VGND VGND VPWR VPWR _17871_/C sky130_fd_sc_hd__nand2_4
XFILLER_61_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16821_ _14913_/Y _16819_/X HWDATA[18] _16819_/X VGND VGND VPWR VPWR _24419_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15184__B _15165_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19928__B1 _19841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16752_ _24452_/Q VGND VGND VPWR VPWR _16752_/Y sky130_fd_sc_hd__inv_2
X_19540_ _19534_/Y _19539_/X _19426_/X _19539_/X VGND VGND VPWR VPWR _19540_/X sky130_fd_sc_hd__a2bb2o_4
X_13964_ _13931_/Y _13964_/B _13950_/X _13963_/X VGND VGND VPWR VPWR _13964_/X sky130_fd_sc_hd__or4_4
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15703_ _15703_/A VGND VGND VPWR VPWR _15742_/A sky130_fd_sc_hd__inv_2
X_12915_ _12753_/X _12903_/X VGND VGND VPWR VPWR _12915_/X sky130_fd_sc_hd__or2_4
XANTENNA__18600__B1 _16541_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16683_ _16664_/A VGND VGND VPWR VPWR _16683_/X sky130_fd_sc_hd__buf_2
X_19471_ _19470_/Y VGND VGND VPWR VPWR _19471_/X sky130_fd_sc_hd__buf_2
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13895_ _13895_/A VGND VGND VPWR VPWR _13895_/X sky130_fd_sc_hd__buf_2
XFILLER_34_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16296__A _16288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15634_ _24882_/Q VGND VGND VPWR VPWR _21584_/A sky130_fd_sc_hd__inv_2
X_18422_ _18422_/A _18417_/X _18419_/X _18422_/D VGND VGND VPWR VPWR _18422_/X sky130_fd_sc_hd__or4_4
X_12846_ _12955_/A _12846_/B _12944_/C _12941_/A VGND VGND VPWR VPWR _12846_/X sky130_fd_sc_hd__or4_4
XFILLER_61_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18353_ _18350_/Y _17478_/X _18352_/Y VGND VGND VPWR VPWR _18353_/Y sky130_fd_sc_hd__o21ai_4
X_15565_ _15565_/A VGND VGND VPWR VPWR _15565_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_247_0_HCLK clkbuf_8_247_0_HCLK/A VGND VGND VPWR VPWR _25024_/CLK sky130_fd_sc_hd__clkbuf_1
X_12777_ _12766_/X _12777_/B _12773_/X _12777_/D VGND VGND VPWR VPWR _12791_/C sky130_fd_sc_hd__or4_4
XPHY_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23977__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17304_ _17279_/A _17304_/B _17303_/X VGND VGND VPWR VPWR _17305_/A sky130_fd_sc_hd__or3_4
XANTENNA__22745__B _23035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _25096_/Q _14511_/X _25095_/Q _14513_/X VGND VGND VPWR VPWR _14516_/X sky130_fd_sc_hd__o22a_4
XPHY_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _11728_/A _11728_/B VGND VGND VPWR VPWR _11730_/C sky130_fd_sc_hd__or2_4
X_18284_ _18275_/X _18278_/X _19930_/A VGND VGND VPWR VPWR _18284_/X sky130_fd_sc_hd__o21a_4
X_15496_ _12050_/X _15494_/X HADDR[21] _15494_/X VGND VGND VPWR VPWR _15496_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20546__A _14381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12571__A2_N _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17235_ _24358_/Q VGND VGND VPWR VPWR _17235_/Y sky130_fd_sc_hd__inv_2
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14447_ _14446_/Y _14442_/X _14403_/X _14442_/X VGND VGND VPWR VPWR _25120_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11659_ _13693_/A VGND VGND VPWR VPWR _11659_/Y sky130_fd_sc_hd__inv_2
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17166_ _16336_/Y _17240_/A _16336_/Y _17240_/A VGND VGND VPWR VPWR _17172_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20069__A3 _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14378_ _14378_/A VGND VGND VPWR VPWR _18895_/A sky130_fd_sc_hd__buf_2
XFILLER_31_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22761__A _23097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16117_ _22902_/A VGND VGND VPWR VPWR _16117_/Y sky130_fd_sc_hd__inv_2
X_13329_ _13426_/A _23617_/Q VGND VGND VPWR VPWR _13329_/X sky130_fd_sc_hd__or2_4
X_17097_ _17108_/A _17095_/X _17096_/X VGND VGND VPWR VPWR _24381_/D sky130_fd_sc_hd__and3_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16048_ _16046_/Y _16047_/X _11818_/X _16047_/X VGND VGND VPWR VPWR _16048_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24765__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19807_ _19807_/A VGND VGND VPWR VPWR _19807_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17999_ _17999_/A _23867_/Q VGND VGND VPWR VPWR _18000_/C sky130_fd_sc_hd__or2_4
XFILLER_84_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19919__B1 _19787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17590__A _17885_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19738_ _19737_/Y _19735_/X _19715_/X _19735_/X VGND VGND VPWR VPWR _23625_/D sky130_fd_sc_hd__a2bb2o_4
X_19669_ _19676_/A VGND VGND VPWR VPWR _19669_/X sky130_fd_sc_hd__buf_2
XFILLER_64_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_57_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21700_ _21108_/B VGND VGND VPWR VPWR _21700_/X sky130_fd_sc_hd__buf_2
XFILLER_53_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22680_ _22671_/A _22669_/Y _22671_/Y _22675_/Y _22679_/Y VGND VGND VPWR VPWR _22680_/X
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__22936__A _24554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21631_ _21631_/A _21631_/B _21631_/C VGND VGND VPWR VPWR _21631_/X sky130_fd_sc_hd__and3_4
XANTENNA__22151__B1 _22885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22655__B _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24350_ _24355_/CLK _17305_/Y HRESETn VGND VGND VPWR VPWR _23008_/A sky130_fd_sc_hd__dfrtp_4
X_21562_ _16453_/B VGND VGND VPWR VPWR _21562_/X sky130_fd_sc_hd__buf_2
XFILLER_138_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13719__B1 _13714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23301_ _24766_/Q _23269_/B VGND VGND VPWR VPWR _23301_/X sky130_fd_sc_hd__or2_4
X_20513_ _20458_/D _20458_/B _20513_/C _20513_/D VGND VGND VPWR VPWR _20513_/X sky130_fd_sc_hd__or4_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21493_ _21821_/A VGND VGND VPWR VPWR _21493_/X sky130_fd_sc_hd__buf_2
X_24281_ _24278_/CLK _17692_/X HRESETn VGND VGND VPWR VPWR _17573_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20444_ _20444_/A _20439_/X VGND VGND VPWR VPWR _20453_/A sky130_fd_sc_hd__and2_4
XFILLER_88_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23232_ _23232_/A _23057_/X VGND VGND VPWR VPWR _23235_/B sky130_fd_sc_hd__or2_4
XFILLER_88_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22671__A _22671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17765__A _16916_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20375_ _23389_/Q VGND VGND VPWR VPWR _20375_/Y sky130_fd_sc_hd__inv_2
X_23163_ _20790_/Y _22988_/X _20929_/Y _22790_/X VGND VGND VPWR VPWR _23163_/X sky130_fd_sc_hd__o22a_4
XFILLER_49_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22390__B _22390_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22114_ _14263_/Y _21548_/B _17423_/Y _21549_/B VGND VGND VPWR VPWR _22114_/X sky130_fd_sc_hd__o22a_4
X_23094_ _23071_/X _23075_/X _23094_/C _23094_/D VGND VGND VPWR VPWR HRDATA[24] sky130_fd_sc_hd__or4_4
XFILLER_0_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22045_ _22575_/A VGND VGND VPWR VPWR _22506_/B sky130_fd_sc_hd__buf_2
XANTENNA__15285__A _15165_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21965__B1 _13784_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14620__C _13598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18830__B1 _16539_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24435__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21734__B _22695_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21717__B1 _15473_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23996_ _23995_/CLK _20499_/X HRESETn VGND VGND VPWR VPWR _23996_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22947_ _21409_/A _22945_/X _22826_/X _22946_/X VGND VGND VPWR VPWR _22948_/A sky130_fd_sc_hd__o22a_4
XFILLER_28_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12700_ _12699_/X VGND VGND VPWR VPWR _12700_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13680_ _13721_/A VGND VGND VPWR VPWR _13680_/X sky130_fd_sc_hd__buf_2
XFILLER_70_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22878_ _22878_/A _22796_/B VGND VGND VPWR VPWR _22882_/B sky130_fd_sc_hd__or2_4
XANTENNA__22846__A _22836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12631_ _12625_/B _12631_/B _12631_/C VGND VGND VPWR VPWR _12632_/A sky130_fd_sc_hd__or3_4
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24617_ _24346_/CLK _24617_/D HRESETn VGND VGND VPWR VPWR _22860_/A sky130_fd_sc_hd__dfrtp_4
X_21829_ _21829_/A VGND VGND VPWR VPWR _21829_/Y sky130_fd_sc_hd__inv_2
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22142__B1 _12345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ _15285_/X VGND VGND VPWR VPWR _15372_/A sky130_fd_sc_hd__buf_2
XANTENNA__25294__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_0_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12562_ _12562_/A VGND VGND VPWR VPWR _12562_/Y sky130_fd_sc_hd__inv_2
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24548_ _24517_/CLK _24548_/D HRESETn VGND VGND VPWR VPWR _16503_/A sky130_fd_sc_hd__dfrtp_4
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_14_0_HCLK clkbuf_7_7_0_HCLK/X VGND VGND VPWR VPWR _23581_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14301_ _13643_/B _14301_/B _14300_/X VGND VGND VPWR VPWR _25167_/D sky130_fd_sc_hd__and3_4
XANTENNA__22780__A1_N _17253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25223__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15281_ _15278_/A _15278_/B VGND VGND VPWR VPWR _15281_/Y sky130_fd_sc_hd__nand2_4
XFILLER_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _12471_/D VGND VGND VPWR VPWR _12494_/B sky130_fd_sc_hd__inv_2
Xclkbuf_8_77_0_HCLK clkbuf_8_77_0_HCLK/A VGND VGND VPWR VPWR _24942_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24479_ _24496_/CLK _24479_/D HRESETn VGND VGND VPWR VPWR _24479_/Q sky130_fd_sc_hd__dfrtp_4
X_17020_ _17260_/A VGND VGND VPWR VPWR _17020_/X sky130_fd_sc_hd__buf_2
XFILLER_32_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ _14231_/Y _14229_/X _13797_/X _14229_/X VGND VGND VPWR VPWR _14232_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22445__A1 _16518_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18649__B1 _24523_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22445__B2 _16795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14163_ _14129_/X _14162_/X _25121_/Q _14132_/A VGND VGND VPWR VPWR _14163_/Y sky130_fd_sc_hd__a22oi_4
X_13114_ _25323_/Q _13114_/B VGND VGND VPWR VPWR _13115_/B sky130_fd_sc_hd__or2_4
XANTENNA__21197__A _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14094_ _14394_/A VGND VGND VPWR VPWR _14381_/A sky130_fd_sc_hd__inv_2
X_18971_ _23890_/Q VGND VGND VPWR VPWR _18971_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20208__B1 _20123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15883__B1 _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21405__C1 _21404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13045_ _12990_/B _13045_/B VGND VGND VPWR VPWR _13048_/B sky130_fd_sc_hd__or2_4
X_17922_ _13541_/C _17921_/Y _17916_/X VGND VGND VPWR VPWR _17922_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19074__B1 _18977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17853_ _17744_/A _17853_/B VGND VGND VPWR VPWR _17855_/B sky130_fd_sc_hd__or2_4
XANTENNA__15635__B1 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16804_ _14967_/Y _16802_/X HWDATA[28] _16802_/X VGND VGND VPWR VPWR _24429_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24105__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14996_ _14996_/A _14996_/B _14992_/X _14996_/D VGND VGND VPWR VPWR _15022_/A sky130_fd_sc_hd__or4_4
X_17784_ _17786_/B VGND VGND VPWR VPWR _17790_/B sky130_fd_sc_hd__inv_2
XFILLER_47_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23173__A2 _22998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19523_ _19523_/A VGND VGND VPWR VPWR _19523_/Y sky130_fd_sc_hd__inv_2
X_13947_ _13947_/A _13947_/B VGND VGND VPWR VPWR _13950_/C sky130_fd_sc_hd__nor2_4
X_16735_ _15005_/Y _16730_/X _16380_/X _16734_/X VGND VGND VPWR VPWR _16735_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16666_ _24488_/Q VGND VGND VPWR VPWR _16666_/Y sky130_fd_sc_hd__inv_2
X_19454_ _18073_/B VGND VGND VPWR VPWR _19454_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13878_ _25233_/Q _13860_/X _25232_/Q _13855_/X VGND VGND VPWR VPWR _13878_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14258__B _14223_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15617_ _15561_/X VGND VGND VPWR VPWR _15617_/X sky130_fd_sc_hd__buf_2
X_18405_ _24164_/Q VGND VGND VPWR VPWR _18405_/Y sky130_fd_sc_hd__inv_2
X_12829_ _12845_/A _24775_/Q _25356_/Q _12795_/Y VGND VGND VPWR VPWR _12829_/X sky130_fd_sc_hd__a2bb2o_4
X_16597_ _16597_/A VGND VGND VPWR VPWR _16597_/Y sky130_fd_sc_hd__inv_2
X_19385_ _19383_/Y _19379_/X _19294_/X _19384_/X VGND VGND VPWR VPWR _23746_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15548_ _15728_/A VGND VGND VPWR VPWR _15548_/X sky130_fd_sc_hd__buf_2
X_18336_ _18333_/X _18335_/X _18333_/X _18335_/X VGND VGND VPWR VPWR _18336_/X sky130_fd_sc_hd__a2bb2o_4
X_18267_ HWDATA[1] VGND VGND VPWR VPWR _18267_/X sky130_fd_sc_hd__buf_2
X_15479_ _14876_/Y _15476_/X _14470_/X _15476_/X VGND VGND VPWR VPWR _24939_/D sky130_fd_sc_hd__a2bb2o_4
X_17218_ _24356_/Q VGND VGND VPWR VPWR _17234_/A sky130_fd_sc_hd__inv_2
X_18198_ _17995_/A _18198_/B _18198_/C VGND VGND VPWR VPWR _18198_/X sky130_fd_sc_hd__and3_4
XFILLER_11_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17149_ _17130_/B VGND VGND VPWR VPWR _17149_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24946__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20160_ _20160_/A VGND VGND VPWR VPWR _21616_/B sky130_fd_sc_hd__inv_2
XFILLER_89_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21538__C _21095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20091_ _23496_/Q VGND VGND VPWR VPWR _20091_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21947__B1 _18298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23850_ _24396_/CLK _19092_/X VGND VGND VPWR VPWR _19090_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22801_ _23021_/A _22801_/B _22801_/C VGND VGND VPWR VPWR _22806_/C sky130_fd_sc_hd__and3_4
XFILLER_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23781_ _23846_/CLK _19283_/X VGND VGND VPWR VPWR _23781_/Q sky130_fd_sc_hd__dfxtp_4
X_20993_ _20992_/A _20992_/B _24326_/Q _20992_/X VGND VGND VPWR VPWR _23966_/D sky130_fd_sc_hd__o22a_4
X_25520_ _24275_/CLK _11810_/X HRESETn VGND VGND VPWR VPWR _25520_/Q sky130_fd_sc_hd__dfrtp_4
X_22732_ _22731_/X VGND VGND VPWR VPWR _22732_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15929__A1 _15669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22666__A _16506_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21570__A _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25182__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25451_ _25368_/CLK _12389_/X HRESETn VGND VGND VPWR VPWR _25451_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22663_ _22662_/X VGND VGND VPWR VPWR _22663_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16664__A _16664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24402_ _24596_/CLK _24402_/D HRESETn VGND VGND VPWR VPWR _14944_/A sky130_fd_sc_hd__dfrtp_4
X_21614_ _21614_/A _21606_/X _21613_/X VGND VGND VPWR VPWR _21614_/X sky130_fd_sc_hd__or3_4
X_25382_ _25356_/CLK _25382_/D HRESETn VGND VGND VPWR VPWR _12747_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_230_0_HCLK clkbuf_8_230_0_HCLK/A VGND VGND VPWR VPWR _24830_/CLK sky130_fd_sc_hd__clkbuf_1
X_22594_ _21064_/A _22591_/X _21098_/X _22593_/X VGND VGND VPWR VPWR _22594_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_90_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24333_ _24177_/CLK _17373_/X HRESETn VGND VGND VPWR VPWR _24333_/Q sky130_fd_sc_hd__dfrtp_4
X_21545_ _21540_/X _21542_/Y _21543_/X _21544_/X VGND VGND VPWR VPWR _21545_/X sky130_fd_sc_hd__and4_4
XFILLER_138_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22427__B2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24264_ _24689_/CLK _17820_/X HRESETn VGND VGND VPWR VPWR _24264_/Q sky130_fd_sc_hd__dfrtp_4
X_21476_ _21454_/A VGND VGND VPWR VPWR _21485_/A sky130_fd_sc_hd__buf_2
XFILLER_14_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23215_ _23274_/A _23214_/X VGND VGND VPWR VPWR _23222_/C sky130_fd_sc_hd__and2_4
X_20427_ _20445_/B _20444_/A _20427_/C VGND VGND VPWR VPWR _20428_/D sky130_fd_sc_hd__or3_4
XANTENNA__24687__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24195_ _24186_/CLK _18336_/X HRESETn VGND VGND VPWR VPWR _24195_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23146_ _23274_/A _23145_/X VGND VGND VPWR VPWR _23155_/C sky130_fd_sc_hd__and2_4
X_20358_ _20358_/A VGND VGND VPWR VPWR _22346_/B sky130_fd_sc_hd__inv_2
XANTENNA__24616__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20289_ _23422_/Q VGND VGND VPWR VPWR _20289_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_2_0_HCLK_A clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23077_ _12277_/B _22820_/X _23076_/X VGND VGND VPWR VPWR _23077_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_114_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22028_ _22005_/X _22028_/B VGND VGND VPWR VPWR _22028_/X sky130_fd_sc_hd__or2_4
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14850_ _14828_/X _14849_/X _25181_/Q _14835_/X VGND VGND VPWR VPWR _14850_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_114_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15743__A HWDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13801_ _13799_/Y _13796_/X _13800_/X _13796_/X VGND VGND VPWR VPWR _25261_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16290__B1 _15940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14781_ _14781_/A _14781_/B VGND VGND VPWR VPWR _14781_/X sky130_fd_sc_hd__and2_4
XANTENNA__15462__B _14223_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11993_ _24088_/Q _11992_/X VGND VGND VPWR VPWR _11994_/B sky130_fd_sc_hd__and2_4
XFILLER_21_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23979_ _25219_/CLK _23979_/D HRESETn VGND VGND VPWR VPWR _20650_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16520_ _24541_/Q VGND VGND VPWR VPWR _16520_/Y sky130_fd_sc_hd__inv_2
X_13732_ _13729_/B _13731_/X _13680_/X _13714_/A _11682_/A VGND VGND VPWR VPWR _25269_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25475__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_40_0_HCLK clkbuf_6_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_81_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16451_ _16451_/A VGND VGND VPWR VPWR _16452_/A sky130_fd_sc_hd__buf_2
XANTENNA__25404__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13663_ _13663_/A _13663_/B _24044_/Q _20879_/A VGND VGND VPWR VPWR _20900_/A sky130_fd_sc_hd__or4_4
XFILLER_95_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15402_ _15299_/B _15392_/X VGND VGND VPWR VPWR _15403_/C sky130_fd_sc_hd__nand2_4
X_12614_ _12731_/A _12729_/A _12510_/Y _12712_/A VGND VGND VPWR VPWR _12614_/X sky130_fd_sc_hd__or4_4
X_19170_ _19169_/Y _19167_/X _19056_/X _19167_/X VGND VGND VPWR VPWR _23822_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16382_ _16389_/A VGND VGND VPWR VPWR _16382_/X sky130_fd_sc_hd__buf_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13594_ _24913_/Q _15542_/A VGND VGND VPWR VPWR _13595_/A sky130_fd_sc_hd__or2_4
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18121_ _18185_/A _18121_/B _18120_/X VGND VGND VPWR VPWR _18129_/B sky130_fd_sc_hd__or3_4
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15333_ _15325_/B _15316_/X _15087_/Y VGND VGND VPWR VPWR _15333_/X sky130_fd_sc_hd__o21a_4
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12545_ _25417_/Q VGND VGND VPWR VPWR _12636_/A sky130_fd_sc_hd__inv_2
XANTENNA__21874__C1 _21095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14094__A _14394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18052_ _18187_/A _19159_/A VGND VGND VPWR VPWR _18053_/C sky130_fd_sc_hd__or2_4
X_15264_ _15251_/B _15250_/X _15190_/A _15261_/B VGND VGND VPWR VPWR _15265_/A sky130_fd_sc_hd__a211o_4
X_12476_ _12503_/A _12476_/B _12476_/C VGND VGND VPWR VPWR _12476_/X sky130_fd_sc_hd__and3_4
XFILLER_126_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17003_ _17003_/A _17003_/B _17001_/X _17002_/X VGND VGND VPWR VPWR _17003_/X sky130_fd_sc_hd__or4_4
XFILLER_6_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14215_ _14214_/Y _14210_/X _13810_/X _14201_/A VGND VGND VPWR VPWR _14215_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15195_ _15194_/X VGND VGND VPWR VPWR _15195_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14146_ _14132_/A VGND VGND VPWR VPWR _14146_/X sky130_fd_sc_hd__buf_2
XANTENNA__24357__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14077_ _13998_/X _14065_/X _14057_/X _13997_/X _14076_/X VGND VGND VPWR VPWR _14077_/X
+ sky130_fd_sc_hd__a32o_4
X_18954_ _13308_/B VGND VGND VPWR VPWR _18954_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13028_ _13043_/A _13043_/B _12999_/B _13028_/D VGND VGND VPWR VPWR _13029_/B sky130_fd_sc_hd__or4_4
X_17905_ _17905_/A VGND VGND VPWR VPWR _17905_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18885_ _20562_/A VGND VGND VPWR VPWR _20582_/B sky130_fd_sc_hd__buf_2
XANTENNA__15608__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15653__A _15653_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17836_ _17835_/X VGND VGND VPWR VPWR _24259_/D sky130_fd_sc_hd__inv_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_122_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_245_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17767_ _23314_/A _17768_/B VGND VGND VPWR VPWR _17767_/X sky130_fd_sc_hd__or2_4
X_14979_ _25023_/Q _14967_/Y _15249_/A _24405_/Q VGND VGND VPWR VPWR _14979_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23992__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19506_ _19506_/A VGND VGND VPWR VPWR _19506_/Y sky130_fd_sc_hd__inv_2
X_16718_ _16716_/Y _16712_/X _16717_/X _16712_/X VGND VGND VPWR VPWR _24467_/D sky130_fd_sc_hd__a2bb2o_4
X_17698_ _17577_/Y _17600_/D _17601_/X _17696_/B VGND VGND VPWR VPWR _17699_/A sky130_fd_sc_hd__a211o_4
XFILLER_62_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23921__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24106__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25145__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19437_ _18140_/B VGND VGND VPWR VPWR _19437_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16649_ _16648_/Y _16646_/X _16380_/X _16646_/X VGND VGND VPWR VPWR _24495_/D sky130_fd_sc_hd__a2bb2o_4
X_19368_ _18132_/B VGND VGND VPWR VPWR _19368_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18319_ _17700_/X _18319_/B _18319_/C VGND VGND VPWR VPWR _18319_/X sky130_fd_sc_hd__or3_4
XFILLER_37_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19299_ _19299_/A VGND VGND VPWR VPWR _19299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17533__B1 _11807_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21330_ _14377_/B _21350_/B VGND VGND VPWR VPWR _21331_/A sky130_fd_sc_hd__or2_4
XFILLER_11_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_60_0_HCLK clkbuf_8_61_0_HCLK/A VGND VGND VPWR VPWR _24720_/CLK sky130_fd_sc_hd__clkbuf_1
X_21261_ _21244_/X _21259_/X _21260_/X VGND VGND VPWR VPWR _21261_/X sky130_fd_sc_hd__a21o_4
XANTENNA__24780__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21549__B _21549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23000_ _24422_/Q _22929_/X _22997_/X _22999_/X VGND VGND VPWR VPWR _23000_/X sky130_fd_sc_hd__a211o_4
X_20212_ _20211_/Y VGND VGND VPWR VPWR _20212_/X sky130_fd_sc_hd__buf_2
XFILLER_102_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21192_ _21192_/A _19968_/Y VGND VGND VPWR VPWR _21194_/B sky130_fd_sc_hd__or2_4
XANTENNA__24098__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15847__B1 _12604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20143_ _20142_/Y _20140_/X _20099_/X _20140_/X VGND VGND VPWR VPWR _23478_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24027__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12252__A _12252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20074_ _20065_/A _18325_/X _11862_/A _13412_/B _20065_/Y VGND VGND VPWR VPWR _23502_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_44_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24951_ _24950_/CLK _15454_/X HRESETn VGND VGND VPWR VPWR _13909_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_100_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22593__B1 _24714_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15563__A _15563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23902_ _24209_/CLK _18941_/X VGND VGND VPWR VPWR _13411_/B sky130_fd_sc_hd__dfxtp_4
X_24882_ _24643_/CLK _24882_/D HRESETn VGND VGND VPWR VPWR _24882_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23833_ _25264_/CLK _23833_/D VGND VGND VPWR VPWR _19139_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22345__B1 _21679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23764_ _23828_/CLK _23764_/D VGND VGND VPWR VPWR _17933_/B sky130_fd_sc_hd__dfxtp_4
X_20976_ _20976_/A VGND VGND VPWR VPWR _20978_/A sky130_fd_sc_hd__inv_2
XFILLER_81_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22396__A _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_27_0_HCLK clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_25503_ _25503_/CLK _25503_/D HRESETn VGND VGND VPWR VPWR _11870_/A sky130_fd_sc_hd__dfrtp_4
X_22715_ _24749_/Q _22265_/X _15894_/A _24821_/Q _22426_/X VGND VGND VPWR VPWR _22716_/A
+ sky130_fd_sc_hd__a32o_4
X_23695_ _23711_/CLK _19529_/X VGND VGND VPWR VPWR _19527_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25434_ _25425_/CLK _25434_/D HRESETn VGND VGND VPWR VPWR _25434_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22648__A1 _15709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22646_ _22646_/A _22645_/X VGND VGND VPWR VPWR _22658_/B sky130_fd_sc_hd__and2_4
XANTENNA__22648__B2 _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25365_ _25356_/CLK _25365_/D HRESETn VGND VGND VPWR VPWR _12843_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_16_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24868__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22577_ _11671_/Y _22727_/B VGND VGND VPWR VPWR _22577_/X sky130_fd_sc_hd__and2_4
X_12330_ _12330_/A VGND VGND VPWR VPWR _13092_/A sky130_fd_sc_hd__inv_2
X_24316_ _24883_/CLK _24316_/D HRESETn VGND VGND VPWR VPWR _24316_/Q sky130_fd_sc_hd__dfrtp_4
X_21528_ _21528_/A VGND VGND VPWR VPWR _21528_/Y sky130_fd_sc_hd__inv_2
X_25296_ _25301_/CLK _13513_/X HRESETn VGND VGND VPWR VPWR _25296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12261_ _12252_/A _12259_/Y _12433_/A _12257_/A VGND VGND VPWR VPWR _12261_/X sky130_fd_sc_hd__a2bb2o_4
X_24247_ _24673_/CLK _17882_/X HRESETn VGND VGND VPWR VPWR _24247_/Q sky130_fd_sc_hd__dfrtp_4
X_21459_ _21459_/A _20038_/Y VGND VGND VPWR VPWR _21460_/C sky130_fd_sc_hd__or2_4
XANTENNA__12355__A2_N _24830_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14000_ _25227_/Q VGND VGND VPWR VPWR _14001_/D sky130_fd_sc_hd__buf_2
XFILLER_123_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24450__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12192_ _25430_/Q _12190_/Y _12290_/A _24761_/Q VGND VGND VPWR VPWR _12198_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24178_ _23933_/CLK _18388_/X HRESETn VGND VGND VPWR VPWR _24178_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15838__B1 _24810_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13258__A _13195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23129_ _23129_/A _23057_/X VGND VGND VPWR VPWR _23129_/X sky130_fd_sc_hd__or2_4
XFILLER_62_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15951_ _15930_/X _15935_/X HWDATA[23] _24758_/Q _15933_/X VGND VGND VPWR VPWR _15951_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_27_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22584__B1 _22527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16569__A _24523_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14902_ _25005_/Q _14900_/Y _15071_/A _24427_/Q VGND VGND VPWR VPWR _14910_/B sky130_fd_sc_hd__a2bb2o_4
X_15882_ _15868_/X VGND VGND VPWR VPWR _15882_/X sky130_fd_sc_hd__buf_2
X_18670_ _18742_/A VGND VGND VPWR VPWR _18738_/A sky130_fd_sc_hd__buf_2
XFILLER_114_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17621_ _17581_/X _17600_/D _17543_/Y VGND VGND VPWR VPWR _17621_/X sky130_fd_sc_hd__o21a_4
XFILLER_40_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14833_ _23987_/D _14832_/X _25186_/Q _23987_/D VGND VGND VPWR VPWR _25041_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15192__B _15069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14764_ _14763_/X VGND VGND VPWR VPWR _14764_/Y sky130_fd_sc_hd__inv_2
X_17552_ _17524_/X _17551_/X VGND VGND VPWR VPWR _17792_/C sky130_fd_sc_hd__or2_4
XANTENNA__19201__B1 _19133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11976_ _11976_/A _11975_/X VGND VGND VPWR VPWR _11976_/X sky130_fd_sc_hd__and2_4
XFILLER_17_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13715_ _13689_/X _13707_/X _13712_/Y _13714_/X _25277_/Q VGND VGND VPWR VPWR _25277_/D
+ sky130_fd_sc_hd__a32o_4
X_16503_ _16503_/A VGND VGND VPWR VPWR _16503_/Y sky130_fd_sc_hd__inv_2
X_17483_ _24196_/Q _17468_/X VGND VGND VPWR VPWR _17483_/X sky130_fd_sc_hd__and2_4
X_14695_ _21612_/A _14694_/X _21612_/A _14694_/X VGND VGND VPWR VPWR _14719_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19222_ _19221_/Y VGND VGND VPWR VPWR _19222_/X sky130_fd_sc_hd__buf_2
XFILLER_72_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13646_ _25287_/Q _13644_/X _13673_/A VGND VGND VPWR VPWR _24084_/D sky130_fd_sc_hd__o21ai_4
X_16434_ _15077_/Y _16433_/X _16061_/X _16433_/X VGND VGND VPWR VPWR _24573_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22639__B2 _22429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16365_ _24599_/Q VGND VGND VPWR VPWR _16365_/Y sky130_fd_sc_hd__inv_2
X_19153_ _19153_/A VGND VGND VPWR VPWR _19153_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13577_ _13575_/A _13576_/A _13575_/Y _13576_/Y VGND VGND VPWR VPWR _13578_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12337__A _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15316_ _15310_/B _15165_/B VGND VGND VPWR VPWR _15316_/X sky130_fd_sc_hd__and2_4
X_18104_ _18104_/A _20221_/A VGND VGND VPWR VPWR _18105_/C sky130_fd_sc_hd__or2_4
X_12528_ _25409_/Q _12526_/Y _25415_/Q _12527_/Y VGND VGND VPWR VPWR _12528_/X sky130_fd_sc_hd__a2bb2o_4
X_16296_ _16288_/X VGND VGND VPWR VPWR _16296_/X sky130_fd_sc_hd__buf_2
X_19084_ _20043_/C _20043_/D _13735_/X _19084_/D VGND VGND VPWR VPWR _19084_/X sky130_fd_sc_hd__or4_4
XANTENNA__24538__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17847__B _17792_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_47_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15247_ _14908_/X _15171_/B VGND VGND VPWR VPWR _15248_/B sky130_fd_sc_hd__or2_4
X_18035_ _18201_/A _18033_/X _18035_/C VGND VGND VPWR VPWR _18039_/B sky130_fd_sc_hd__and3_4
XANTENNA__15648__A _15648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12459_ _12283_/X _13008_/B VGND VGND VPWR VPWR _12459_/X sky130_fd_sc_hd__or2_4
XFILLER_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18024__A _18024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15178_ _15180_/B VGND VGND VPWR VPWR _15179_/B sky130_fd_sc_hd__inv_2
XANTENNA__24191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14129_ _14129_/A VGND VGND VPWR VPWR _14129_/X sky130_fd_sc_hd__buf_2
XANTENNA__20822__B1 _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24120__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19986_ _21938_/B _19982_/X _19985_/X _19982_/X VGND VGND VPWR VPWR _19986_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12072__A _16183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25354__CLK _25354_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18937_ _18937_/A VGND VGND VPWR VPWR _18937_/X sky130_fd_sc_hd__buf_2
XANTENNA__25397__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18868_ _18884_/A VGND VGND VPWR VPWR _18868_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25326__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17819_ _16914_/Y _17824_/B _16955_/X VGND VGND VPWR VPWR _17819_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_67_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18799_ _18799_/A _18797_/X _18798_/X VGND VGND VPWR VPWR _24122_/D sky130_fd_sc_hd__and3_4
X_20830_ _16711_/Y _20815_/X _20824_/X _20829_/X VGND VGND VPWR VPWR _20830_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16006__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23105__A _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20761_ _20761_/A _13120_/D VGND VGND VPWR VPWR _20761_/X sky130_fd_sc_hd__or2_4
XFILLER_39_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22500_ _22671_/A _22500_/B VGND VGND VPWR VPWR _22518_/A sky130_fd_sc_hd__nor2_4
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23480_ _23496_/CLK _23480_/D VGND VGND VPWR VPWR _23480_/Q sky130_fd_sc_hd__dfxtp_4
X_20692_ _21739_/A _20677_/X _20686_/X _20691_/X VGND VGND VPWR VPWR _20692_/X sky130_fd_sc_hd__o22a_4
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22431_ _12769_/Y _21858_/X _22272_/X _12536_/Y _21413_/X VGND VGND VPWR VPWR _22431_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_52_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15780__A2 _15669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24961__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25150_ _24109_/CLK _14350_/X HRESETn VGND VGND VPWR VPWR _14338_/A sky130_fd_sc_hd__dfrtp_4
X_22362_ _21885_/X _22360_/X _22362_/C VGND VGND VPWR VPWR _22362_/X sky130_fd_sc_hd__and3_4
XFILLER_104_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21853__A2 _22406_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24279__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24101_ _24102_/CLK _20966_/X HRESETn VGND VGND VPWR VPWR _12151_/A sky130_fd_sc_hd__dfrtp_4
X_21313_ _21556_/A VGND VGND VPWR VPWR _22997_/A sky130_fd_sc_hd__buf_2
XANTENNA__24208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25081_ _25081_/CLK _14588_/X HRESETn VGND VGND VPWR VPWR _25081_/Q sky130_fd_sc_hd__dfrtp_4
X_22293_ _22293_/A _22293_/B _22293_/C _22293_/D VGND VGND VPWR VPWR HRDATA[6] sky130_fd_sc_hd__or4_4
XFILLER_11_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23055__B2 _21211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24032_ _24033_/CLK _24032_/D HRESETn VGND VGND VPWR VPWR _13655_/A sky130_fd_sc_hd__dfrtp_4
X_21244_ _21388_/A _21244_/B _21243_/X VGND VGND VPWR VPWR _21244_/X sky130_fd_sc_hd__or3_4
XFILLER_85_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_4_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21175_ _21186_/A _21172_/X _21174_/X VGND VGND VPWR VPWR _21175_/X sky130_fd_sc_hd__and3_4
XFILLER_78_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20126_ _19844_/X _19084_/D _19822_/C VGND VGND VPWR VPWR _20127_/A sky130_fd_sc_hd__or3_4
XFILLER_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22566__B1 _12282_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20057_ _20057_/A VGND VGND VPWR VPWR _20057_/X sky130_fd_sc_hd__buf_2
X_24934_ _24248_/CLK _24934_/D HRESETn VGND VGND VPWR VPWR _12052_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_19_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16245__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15048__B2 _15027_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20041__B2 _20036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25067__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24865_ _24865_/CLK _15730_/X HRESETn VGND VGND VPWR VPWR _24865_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22838__B _22832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11830_ _11828_/Y _11826_/X _11829_/X _11826_/X VGND VGND VPWR VPWR _11830_/X sky130_fd_sc_hd__a2bb2o_4
X_23816_ _23832_/CLK _19186_/X VGND VGND VPWR VPWR _23816_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22869__B2 _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24796_ _25385_/CLK _15876_/X HRESETn VGND VGND VPWR VPWR _12772_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ HWDATA[26] VGND VGND VPWR VPWR _11761_/X sky130_fd_sc_hd__buf_2
XPHY_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23747_ _23718_/CLK _19382_/X VGND VGND VPWR VPWR _17969_/B sky130_fd_sc_hd__dfxtp_4
X_20959_ _12024_/X _20958_/B VGND VGND VPWR VPWR _20959_/X sky130_fd_sc_hd__and2_4
XPHY_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _12014_/Y _13498_/X _11829_/X _13498_/X VGND VGND VPWR VPWR _25302_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14480_/A VGND VGND VPWR VPWR _14480_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _13689_/A _22507_/A _13689_/A _22507_/A VGND VGND VPWR VPWR _11699_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23678_ _23398_/CLK _23678_/D VGND VGND VPWR VPWR _19576_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22854__A _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _13199_/Y _13415_/X _13430_/X _25315_/Q _11964_/X VGND VGND VPWR VPWR _13431_/X
+ sky130_fd_sc_hd__o32a_4
X_25417_ _25411_/CLK _25417_/D HRESETn VGND VGND VPWR VPWR _25417_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22629_ _21700_/X _22628_/X _21296_/X _16044_/A _21299_/X VGND VGND VPWR VPWR _22629_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_9_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16852__A _16442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16150_ _16149_/Y _16144_/X _16057_/X _16144_/X VGND VGND VPWR VPWR _24675_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13362_ _13426_/A _13362_/B VGND VGND VPWR VPWR _13362_/X sky130_fd_sc_hd__or2_4
X_25348_ _23370_/CLK _25348_/D HRESETn VGND VGND VPWR VPWR _25348_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24631__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15101_ _24987_/Q VGND VGND VPWR VPWR _15338_/A sky130_fd_sc_hd__inv_2
X_12313_ _12313_/A _12313_/B _12313_/C _12312_/X VGND VGND VPWR VPWR _12313_/X sky130_fd_sc_hd__or4_4
XFILLER_6_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16081_ _16079_/A _15674_/X VGND VGND VPWR VPWR _16081_/X sky130_fd_sc_hd__or2_4
XFILLER_5_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23154__A2_N _23149_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13293_ _13162_/X _13293_/B _13292_/X VGND VGND VPWR VPWR _13293_/X sky130_fd_sc_hd__or3_4
X_25279_ _25279_/CLK _13709_/X HRESETn VGND VGND VPWR VPWR _25279_/Q sky130_fd_sc_hd__dfrtp_4
X_15032_ _15227_/A _15030_/Y _15251_/C _15023_/A VGND VGND VPWR VPWR _15032_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12244_ _25443_/Q VGND VGND VPWR VPWR _12244_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19840_ _23589_/Q VGND VGND VPWR VPWR _21223_/B sky130_fd_sc_hd__inv_2
X_12175_ _25452_/Q VGND VGND VPWR VPWR _14329_/A sky130_fd_sc_hd__inv_2
XANTENNA__16484__B1 _16398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19771_ _15845_/A VGND VGND VPWR VPWR _19771_/X sky130_fd_sc_hd__buf_2
XFILLER_3_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16983_ _16983_/A VGND VGND VPWR VPWR _17038_/A sky130_fd_sc_hd__inv_2
XFILLER_110_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16299__A _24624_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18722_ _18733_/A VGND VGND VPWR VPWR _18724_/A sky130_fd_sc_hd__buf_2
XFILLER_67_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25490__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15934_ _15930_/X _15894_/X _15553_/X _24766_/Q _15933_/X VGND VGND VPWR VPWR _24766_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_77_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16236__B1 _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15039__B2 _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21933__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18653_ _16567_/Y _18658_/A _16597_/A _18608_/X VGND VGND VPWR VPWR _18660_/A sky130_fd_sc_hd__a2bb2o_4
X_15865_ _15850_/X _15857_/X _15553_/X _24803_/Q _15864_/X VGND VGND VPWR VPWR _24803_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_64_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17604_ _17604_/A VGND VGND VPWR VPWR _17604_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15931__A _15931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14816_ _25037_/Q _14816_/B _14802_/A VGND VGND VPWR VPWR _14816_/X sky130_fd_sc_hd__or3_4
X_18584_ _18583_/X VGND VGND VPWR VPWR _18584_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15796_ _15781_/X _15795_/X _15714_/X _24837_/Q _15793_/X VGND VGND VPWR VPWR _24837_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_40_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17535_ _11790_/Y _24295_/Q _11776_/A _17630_/A VGND VGND VPWR VPWR _17537_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11959_ _11958_/X _17445_/C VGND VGND VPWR VPWR _11959_/X sky130_fd_sc_hd__or2_4
X_14747_ _21633_/A _14746_/X _21633_/A _14746_/X VGND VGND VPWR VPWR _14747_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17736__B1 _21686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_10_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_14678_ _14691_/A VGND VGND VPWR VPWR _21247_/A sky130_fd_sc_hd__buf_2
X_17466_ _17465_/X VGND VGND VPWR VPWR _17466_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24719__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19205_ _18094_/B VGND VGND VPWR VPWR _19205_/Y sky130_fd_sc_hd__inv_2
X_13629_ _13630_/A VGND VGND VPWR VPWR _18079_/A sky130_fd_sc_hd__inv_2
X_16417_ _16416_/Y _16414_/X _16228_/X _16414_/X VGND VGND VPWR VPWR _16417_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17397_ _20650_/A _20650_/B VGND VGND VPWR VPWR _17398_/B sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_5_5_0_HCLK_A clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19136_ _18996_/X VGND VGND VPWR VPWR _19136_/X sky130_fd_sc_hd__buf_2
X_16348_ _16347_/Y _16343_/X _16057_/X _16343_/X VGND VGND VPWR VPWR _16348_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24372__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12800__A2_N _22623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16279_ _22493_/B _15993_/Y VGND VGND VPWR VPWR _16280_/A sky130_fd_sc_hd__and2_4
X_19067_ _19067_/A VGND VGND VPWR VPWR _19067_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24301__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18018_ _18059_/A _18006_/X _18017_/X VGND VGND VPWR VPWR _18018_/X sky130_fd_sc_hd__and3_4
XFILLER_133_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23499__CLK _23498_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_134_0_HCLK clkbuf_7_67_0_HCLK/X VGND VGND VPWR VPWR _23441_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_102_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16475__B1 _16297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_197_0_HCLK clkbuf_7_98_0_HCLK/X VGND VGND VPWR VPWR _24041_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__25507__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19969_ _19968_/Y _19964_/X _19885_/X _19964_/A VGND VGND VPWR VPWR _19969_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22548__B1 _24852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19413__B1 _19389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22980_ _22714_/A VGND VGND VPWR VPWR _22980_/X sky130_fd_sc_hd__buf_2
XANTENNA__16002__A _15995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21931_ _21912_/X _21929_/X _21930_/X VGND VGND VPWR VPWR _21931_/X sky130_fd_sc_hd__and3_4
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24650_ _24581_/CLK _16226_/X HRESETn VGND VGND VPWR VPWR _16223_/A sky130_fd_sc_hd__dfrtp_4
X_21862_ _21862_/A _21862_/B _21862_/C _21861_/X VGND VGND VPWR VPWR _21862_/X sky130_fd_sc_hd__or4_4
XFILLER_55_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23601_ _23683_/CLK _19811_/X VGND VGND VPWR VPWR _13330_/B sky130_fd_sc_hd__dfxtp_4
X_20813_ _20812_/Y _13668_/X VGND VGND VPWR VPWR _20863_/A sky130_fd_sc_hd__or2_4
XFILLER_36_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24581_ _24581_/CLK _16420_/X HRESETn VGND VGND VPWR VPWR _24581_/Q sky130_fd_sc_hd__dfrtp_4
X_21793_ _21459_/A _21793_/B VGND VGND VPWR VPWR _21794_/C sky130_fd_sc_hd__or2_4
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23532_ _23394_/CLK _20003_/X VGND VGND VPWR VPWR _19999_/A sky130_fd_sc_hd__dfxtp_4
X_20744_ _20761_/A VGND VGND VPWR VPWR _20772_/C sky130_fd_sc_hd__buf_2
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23463_ _24089_/CLK _20183_/X VGND VGND VPWR VPWR _20181_/A sky130_fd_sc_hd__dfxtp_4
X_20675_ _20674_/Y _20675_/B VGND VGND VPWR VPWR _20724_/A sky130_fd_sc_hd__or2_4
XANTENNA__15753__A2 _15742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23276__B2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25202_ _25199_/CLK _25202_/D HRESETn VGND VGND VPWR VPWR _14099_/C sky130_fd_sc_hd__dfrtp_4
X_22414_ _20846_/Y _22278_/X _13129_/A _21304_/X VGND VGND VPWR VPWR _22414_/X sky130_fd_sc_hd__a2bb2o_4
X_23394_ _23394_/CLK _23394_/D VGND VGND VPWR VPWR _23394_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11775__B1 _11774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15288__A _15246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25133_ _25137_/CLK _25133_/D HRESETn VGND VGND VPWR VPWR _20596_/A sky130_fd_sc_hd__dfrtp_4
X_22345_ _22341_/X _22344_/X _21679_/X VGND VGND VPWR VPWR _22345_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24042__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14192__A _14192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23001__C _23000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21039__B1 _22664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_30_0_HCLK clkbuf_7_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_61_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14713__B1 _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25064_ _23826_/CLK _14644_/X HRESETn VGND VGND VPWR VPWR _14785_/A sky130_fd_sc_hd__dfrtp_4
X_22276_ _22658_/A _22276_/B VGND VGND VPWR VPWR _22293_/C sky130_fd_sc_hd__nor2_4
XFILLER_105_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_93_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_93_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_24015_ _24868_/CLK _20760_/X HRESETn VGND VGND VPWR VPWR _13119_/B sky130_fd_sc_hd__dfrtp_4
X_21227_ _14691_/A VGND VGND VPWR VPWR _21377_/A sky130_fd_sc_hd__inv_2
XFILLER_105_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23930__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25248__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21158_ _16445_/Y _21556_/A _16722_/A _21157_/X VGND VGND VPWR VPWR _21158_/X sky130_fd_sc_hd__a211o_4
X_20109_ _22209_/B _20106_/X _20082_/X _20106_/X VGND VGND VPWR VPWR _20109_/X sky130_fd_sc_hd__a2bb2o_4
X_13980_ _13980_/A VGND VGND VPWR VPWR _13980_/Y sky130_fd_sc_hd__inv_2
X_21089_ _21089_/A VGND VGND VPWR VPWR _21089_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12440__A _12199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16218__B1 _15959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12931_ _12602_/A _12847_/X VGND VGND VPWR VPWR _12931_/X sky130_fd_sc_hd__or2_4
XANTENNA__22554__A3 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24917_ _25255_/CLK _15534_/X HRESETn VGND VGND VPWR VPWR _13787_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_111_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16847__A _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12862_ _12600_/X _12838_/A VGND VGND VPWR VPWR _12862_/X sky130_fd_sc_hd__and2_4
X_15650_ _16640_/B _15843_/A VGND VGND VPWR VPWR _15650_/X sky130_fd_sc_hd__or2_4
X_24848_ _23370_/CLK _24848_/D HRESETn VGND VGND VPWR VPWR _12514_/A sky130_fd_sc_hd__dfrtp_4
X_11813_ _11812_/X VGND VGND VPWR VPWR _11813_/X sky130_fd_sc_hd__buf_2
X_14601_ _13559_/Y _14601_/B VGND VGND VPWR VPWR _14601_/Y sky130_fd_sc_hd__nand2_4
X_15581_ _15588_/A VGND VGND VPWR VPWR _15581_/X sky130_fd_sc_hd__buf_2
XFILLER_73_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12793_ _25360_/Q VGND VGND VPWR VPWR _12959_/A sky130_fd_sc_hd__inv_2
XANTENNA__24883__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24779_ _24813_/CLK _15902_/X HRESETn VGND VGND VPWR VPWR _24779_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _21119_/A _14510_/X _23379_/Q _14505_/X VGND VGND VPWR VPWR _14532_/X sky130_fd_sc_hd__o22a_4
X_17320_ _17253_/Y _17320_/B VGND VGND VPWR VPWR _17321_/B sky130_fd_sc_hd__or2_4
XPHY_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11706_/Y _11742_/X _11743_/X _11742_/X VGND VGND VPWR VPWR _11744_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24812__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _25112_/Q VGND VGND VPWR VPWR _14463_/Y sky130_fd_sc_hd__inv_2
X_17251_ _22702_/A VGND VGND VPWR VPWR _17252_/B sky130_fd_sc_hd__inv_2
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _11668_/X _11670_/X _11675_/C _11675_/D VGND VGND VPWR VPWR _11700_/B sky130_fd_sc_hd__or4_4
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15744__A2 _15742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ _13162_/A _13410_/X _13414_/C VGND VGND VPWR VPWR _13415_/C sky130_fd_sc_hd__or3_4
X_16202_ _23129_/A VGND VGND VPWR VPWR _16202_/Y sky130_fd_sc_hd__inv_2
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17182_ _24346_/Q VGND VGND VPWR VPWR _17254_/A sky130_fd_sc_hd__inv_2
XFILLER_122_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14394_ _14394_/A _14394_/B VGND VGND VPWR VPWR _14394_/X sky130_fd_sc_hd__or2_4
XFILLER_128_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16133_ _22655_/A VGND VGND VPWR VPWR _16133_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13345_ _13345_/A _18957_/A VGND VGND VPWR VPWR _13345_/X sky130_fd_sc_hd__or2_4
XFILLER_115_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16064_ _16528_/A VGND VGND VPWR VPWR _16064_/X sky130_fd_sc_hd__buf_2
X_13276_ _13143_/X _13268_/X _13276_/C VGND VGND VPWR VPWR _13276_/X sky130_fd_sc_hd__and3_4
X_15015_ _15015_/A VGND VGND VPWR VPWR _15015_/Y sky130_fd_sc_hd__inv_2
X_12227_ _12186_/X _12198_/X _12212_/X _12227_/D VGND VGND VPWR VPWR _12273_/A sky130_fd_sc_hd__or4_4
XFILLER_68_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_207_0_HCLK clkbuf_8_207_0_HCLK/A VGND VGND VPWR VPWR _24842_/CLK sky130_fd_sc_hd__clkbuf_1
X_19823_ _19823_/A VGND VGND VPWR VPWR _19836_/A sky130_fd_sc_hd__inv_2
X_12158_ _12157_/X VGND VGND VPWR VPWR _20965_/B sky130_fd_sc_hd__buf_2
XFILLER_69_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13446__A _13162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19754_ _13251_/B VGND VGND VPWR VPWR _19754_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12089_ _12088_/Y _12086_/X _11862_/X _12086_/X VGND VGND VPWR VPWR _25467_/D sky130_fd_sc_hd__a2bb2o_4
X_16966_ _24713_/Q _17041_/D _16009_/Y _17026_/A VGND VGND VPWR VPWR _16966_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22759__A _21108_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18705_ _18705_/A _18705_/B _18704_/X VGND VGND VPWR VPWR _18705_/X sky130_fd_sc_hd__or3_4
X_15917_ _15916_/X VGND VGND VPWR VPWR _15917_/Y sky130_fd_sc_hd__inv_2
X_19685_ _19697_/A VGND VGND VPWR VPWR _19685_/X sky130_fd_sc_hd__buf_2
X_16897_ _24255_/Q VGND VGND VPWR VPWR _16898_/A sky130_fd_sc_hd__inv_2
XANTENNA__22478__B _22626_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18636_ _18605_/X _18616_/X _18636_/C _18636_/D VGND VGND VPWR VPWR _18668_/A sky130_fd_sc_hd__or4_4
XANTENNA__19133__A _19642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15848_ _15674_/X _15703_/A VGND VGND VPWR VPWR _15848_/X sky130_fd_sc_hd__or2_4
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23046__A2_N _23042_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18567_ _18471_/Y _18566_/X _18487_/X VGND VGND VPWR VPWR _18567_/Y sky130_fd_sc_hd__a21oi_4
X_15779_ _15777_/A _15674_/X VGND VGND VPWR VPWR _15779_/X sky130_fd_sc_hd__or2_4
XANTENNA__21505__A1 _18272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17518_ _11824_/A _17517_/A _11824_/Y _17517_/Y VGND VGND VPWR VPWR _17518_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24553__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18498_ _18821_/B VGND VGND VPWR VPWR _18498_/X sky130_fd_sc_hd__buf_2
X_17449_ _24310_/Q _17700_/C _17448_/X VGND VGND VPWR VPWR _17449_/X sky130_fd_sc_hd__or3_4
XFILLER_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20460_ _20437_/C _20459_/X VGND VGND VPWR VPWR _20460_/X sky130_fd_sc_hd__or2_4
X_19119_ _19119_/A VGND VGND VPWR VPWR _19119_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20391_ _20383_/X _20379_/X _20072_/X _23382_/Q _20381_/X VGND VGND VPWR VPWR _23382_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22130_ _21589_/X _22128_/X _22130_/C VGND VGND VPWR VPWR _22130_/X sky130_fd_sc_hd__and3_4
XANTENNA__16696__B1 _16340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_17_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22061_ _21885_/X _22059_/X _22060_/X VGND VGND VPWR VPWR _22061_/X sky130_fd_sc_hd__and3_4
XANTENNA__15836__A _15766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21012_ _22764_/A VGND VGND VPWR VPWR _22549_/A sky130_fd_sc_hd__buf_2
XFILLER_138_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21441__B1 _12280_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25341__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16999__B2 _17036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17770__B _17837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22963_ _22963_/A VGND VGND VPWR VPWR _23143_/A sky130_fd_sc_hd__buf_2
XANTENNA__22941__B1 _21050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21914_ _18307_/X VGND VGND VPWR VPWR _21942_/A sky130_fd_sc_hd__buf_2
X_24702_ _24026_/CLK _24702_/D HRESETn VGND VGND VPWR VPWR _21053_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_3_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22894_ _22763_/A _22894_/B VGND VGND VPWR VPWR _22905_/B sky130_fd_sc_hd__and2_4
X_24633_ _24893_/CLK _16272_/X HRESETn VGND VGND VPWR VPWR _21003_/A sky130_fd_sc_hd__dfrtp_4
X_21845_ _21840_/X _21841_/Y _21842_/X _21845_/D VGND VGND VPWR VPWR _21845_/X sky130_fd_sc_hd__and4_4
XFILLER_55_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24294__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24564_ _24561_/CLK _16464_/X HRESETn VGND VGND VPWR VPWR _24564_/Q sky130_fd_sc_hd__dfrtp_4
X_21776_ _14716_/A _21768_/X _21775_/X VGND VGND VPWR VPWR _21776_/X sky130_fd_sc_hd__or3_4
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23515_ _23516_/CLK _20048_/X VGND VGND VPWR VPWR _20047_/A sky130_fd_sc_hd__dfxtp_4
X_20727_ _20721_/X _20723_/Y _15611_/A _20726_/X VGND VGND VPWR VPWR _20727_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24223__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24495_ _24492_/CLK _24495_/D HRESETn VGND VGND VPWR VPWR _16648_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23446_ _23446_/CLK _23446_/D VGND VGND VPWR VPWR _20226_/A sky130_fd_sc_hd__dfxtp_4
X_20658_ _17399_/A _17399_/B _17401_/A VGND VGND VPWR VPWR _20658_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23377_ _23377_/CLK _23377_/D VGND VGND VPWR VPWR _23377_/Q sky130_fd_sc_hd__dfxtp_4
X_20589_ _14405_/Y _20582_/B _18868_/Y _18882_/Y VGND VGND VPWR VPWR _20589_/X sky130_fd_sc_hd__o22a_4
XFILLER_87_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13130_ _24007_/Q _13130_/B VGND VGND VPWR VPWR _13131_/B sky130_fd_sc_hd__or2_4
XFILLER_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25116_ _25113_/CLK _14455_/X HRESETn VGND VGND VPWR VPWR _14394_/A sky130_fd_sc_hd__dfrtp_4
X_22328_ _21944_/A _22328_/B VGND VGND VPWR VPWR _22330_/B sky130_fd_sc_hd__or2_4
XANTENNA__21680__B1 _21679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25429__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17945__B _17945_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22570__C _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13061_ _13061_/A _13064_/B VGND VGND VPWR VPWR _13062_/C sky130_fd_sc_hd__nand2_4
X_25047_ _23516_/CLK _25047_/D HRESETn VGND VGND VPWR VPWR _14762_/C sky130_fd_sc_hd__dfrtp_4
X_22259_ _22259_/A VGND VGND VPWR VPWR _22259_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22224__A2 _22204_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12012_ _12002_/X _12003_/X _12007_/X _12012_/D VGND VGND VPWR VPWR _12012_/X sky130_fd_sc_hd__or4_4
XFILLER_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25082__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16820_ _14927_/Y _16816_/X HWDATA[19] _16819_/X VGND VGND VPWR VPWR _16820_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25011__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_180_0_HCLK clkbuf_7_90_0_HCLK/X VGND VGND VPWR VPWR _24691_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_48_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23185__B1 _24730_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_37_0_HCLK clkbuf_8_37_0_HCLK/A VGND VGND VPWR VPWR _25055_/CLK sky130_fd_sc_hd__clkbuf_1
X_16751_ _15052_/Y _16749_/X _16403_/X _16749_/X VGND VGND VPWR VPWR _24453_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13963_ _13952_/X _13962_/Y VGND VGND VPWR VPWR _13963_/X sky130_fd_sc_hd__or2_4
XANTENNA__21735__A1 _16616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16577__A _24520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22298__B _22298_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15702_ _15702_/A VGND VGND VPWR VPWR _15703_/A sky130_fd_sc_hd__buf_2
XFILLER_19_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12914_ _12850_/C _12912_/X _12913_/Y VGND VGND VPWR VPWR _25374_/D sky130_fd_sc_hd__o21a_4
X_19470_ _19469_/X VGND VGND VPWR VPWR _19470_/Y sky130_fd_sc_hd__inv_2
X_13894_ _13894_/A VGND VGND VPWR VPWR _13918_/D sky130_fd_sc_hd__inv_2
X_16682_ _16682_/A VGND VGND VPWR VPWR _16682_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18421_ _22878_/A _18420_/A _16219_/Y _18420_/Y VGND VGND VPWR VPWR _18422_/D sky130_fd_sc_hd__o22a_4
XFILLER_34_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12845_ _12845_/A _12845_/B _12976_/A VGND VGND VPWR VPWR _12941_/A sky130_fd_sc_hd__or3_4
X_15633_ _21739_/A _15626_/X _15474_/X _15632_/X VGND VGND VPWR VPWR _15633_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18792__A _18792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18352_ _18365_/A _18365_/B VGND VGND VPWR VPWR _18352_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12832__A1_N _25383_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12776_ _25362_/Q _24779_/Q _12774_/Y _12775_/Y VGND VGND VPWR VPWR _12777_/D sky130_fd_sc_hd__o22a_4
X_15564_ _15559_/Y _15563_/X _11746_/X _15563_/X VGND VGND VPWR VPWR _24910_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17256_/X _17267_/X _17222_/Y VGND VGND VPWR VPWR _17303_/X sky130_fd_sc_hd__o21a_4
XPHY_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11727_/A _11727_/B _15523_/A VGND VGND VPWR VPWR _11731_/C sky130_fd_sc_hd__or3_4
X_14515_ _14502_/X _14514_/X VGND VGND VPWR VPWR _25097_/D sky130_fd_sc_hd__or2_4
XFILLER_30_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _15549_/B _15491_/X HADDR[22] _15494_/X VGND VGND VPWR VPWR _24934_/D sky130_fd_sc_hd__a2bb2o_4
X_18283_ _17730_/X _18280_/X _20276_/C VGND VGND VPWR VPWR _19930_/A sky130_fd_sc_hd__or3_4
XFILLER_30_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20171__B1 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17234_ _17234_/A VGND VGND VPWR VPWR _17261_/B sky130_fd_sc_hd__buf_2
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _11656_/Y _21967_/A _13691_/A _24224_/Q VGND VGND VPWR VPWR _11658_/X sky130_fd_sc_hd__a2bb2o_4
X_14446_ _14446_/A VGND VGND VPWR VPWR _14446_/Y sky130_fd_sc_hd__inv_2
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ _15642_/A _14377_/B VGND VGND VPWR VPWR _14378_/A sky130_fd_sc_hd__or2_4
X_17165_ _17164_/X VGND VGND VPWR VPWR _17165_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19864__B1 _19841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12345__A _12345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23946__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13328_ _13234_/A VGND VGND VPWR VPWR _13426_/A sky130_fd_sc_hd__buf_2
X_16116_ _16115_/Y _16113_/X _15957_/X _16113_/X VGND VGND VPWR VPWR _24688_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21658__A _21658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17096_ _17035_/A _17093_/X VGND VGND VPWR VPWR _17096_/X sky130_fd_sc_hd__or2_4
XFILLER_13_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15656__A _15653_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13259_ _13198_/X _13257_/X _25319_/Q _13258_/X VGND VGND VPWR VPWR _25319_/D sky130_fd_sc_hd__o22a_4
X_16047_ _16060_/A VGND VGND VPWR VPWR _16047_/X sky130_fd_sc_hd__buf_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18032__A _18217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19806_ _19805_/Y _19803_/X _19755_/X _19803_/X VGND VGND VPWR VPWR _19806_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17998_ _17990_/A VGND VGND VPWR VPWR _17999_/A sky130_fd_sc_hd__buf_2
XFILLER_81_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19737_ _13325_/B VGND VGND VPWR VPWR _19737_/Y sky130_fd_sc_hd__inv_2
X_16949_ _23219_/A _16948_/X _16156_/Y _17745_/A VGND VGND VPWR VPWR _16949_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19668_ _19668_/A VGND VGND VPWR VPWR _19668_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24734__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_8_0_HCLK clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__16602__B1 _16600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18619_ _24121_/Q VGND VGND VPWR VPWR _18619_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19599_ _18254_/A VGND VGND VPWR VPWR _19599_/X sky130_fd_sc_hd__buf_2
XANTENNA__22936__B _22810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21630_ _21630_/A _20094_/Y VGND VGND VPWR VPWR _21631_/C sky130_fd_sc_hd__or2_4
XFILLER_21_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21561_ _12096_/X VGND VGND VPWR VPWR _21561_/X sky130_fd_sc_hd__buf_2
XANTENNA__15727__A1_N _12539_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20162__B1 _20096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23300_ _23281_/X _23284_/X _23288_/Y _23299_/X VGND VGND VPWR VPWR HRDATA[30] sky130_fd_sc_hd__a211o_4
X_20512_ _23994_/Q _20512_/B VGND VGND VPWR VPWR _20513_/D sky130_fd_sc_hd__and2_4
XFILLER_18_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24280_ _24278_/CLK _17694_/X HRESETn VGND VGND VPWR VPWR _24280_/Q sky130_fd_sc_hd__dfrtp_4
X_21492_ _21260_/X VGND VGND VPWR VPWR _21821_/A sky130_fd_sc_hd__buf_2
XANTENNA__22952__A _23021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23231_ _23128_/A _23230_/X VGND VGND VPWR VPWR _23231_/Y sky130_fd_sc_hd__nor2_4
X_20443_ _20443_/A _20443_/B _20459_/B _20443_/D VGND VGND VPWR VPWR _20443_/X sky130_fd_sc_hd__and4_4
XFILLER_105_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19855__B1 _19787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16669__B1 _16401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25522__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23162_ _23124_/A _23162_/B VGND VGND VPWR VPWR _23162_/Y sky130_fd_sc_hd__nor2_4
X_20374_ _20372_/Y _20373_/X _19629_/A _20373_/X VGND VGND VPWR VPWR _23390_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22113_ _22112_/X VGND VGND VPWR VPWR _22113_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14470__A _14470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19607__B1 _19420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23093_ _23088_/Y _23092_/Y _22850_/X VGND VGND VPWR VPWR _23094_/D sky130_fd_sc_hd__o21a_4
X_22044_ _21504_/B _22044_/B VGND VGND VPWR VPWR _22044_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21965__A1 _21816_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14620__D _14620_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_253_0_HCLK clkbuf_7_126_0_HCLK/X VGND VGND VPWR VPWR _25020_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__13104__C1 _13031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16841__B1 _16600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23995_ _23995_/CLK _20498_/X HRESETn VGND VGND VPWR VPWR _23995_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21717__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13814__A _14406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22946_ _16670_/Y _22790_/A _15587_/Y _22827_/X VGND VGND VPWR VPWR _22946_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24475__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24404__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22877_ _23056_/A _22877_/B VGND VGND VPWR VPWR _22877_/Y sky130_fd_sc_hd__nor2_4
X_12630_ _12623_/C _12629_/X _12623_/A VGND VGND VPWR VPWR _12631_/C sky130_fd_sc_hd__o21a_4
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21828_ _13126_/A _21826_/X _15629_/A _22677_/B VGND VGND VPWR VPWR _21828_/Y sky130_fd_sc_hd__a22oi_4
X_24616_ _24345_/CLK _24616_/D HRESETn VGND VGND VPWR VPWR _22816_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _25405_/Q _12559_/Y _12704_/A _24847_/Q VGND VGND VPWR VPWR _12569_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24547_ _24120_/CLK _16507_/X HRESETn VGND VGND VPWR VPWR _16506_/A sky130_fd_sc_hd__dfrtp_4
X_21759_ _21614_/A _21751_/X _21758_/X VGND VGND VPWR VPWR _21759_/X sky130_fd_sc_hd__or3_4
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14645__A _14645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14300_ _25167_/Q _14299_/Y VGND VGND VPWR VPWR _14300_/X sky130_fd_sc_hd__or2_4
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15280_ _14981_/X _15282_/B _15279_/Y VGND VGND VPWR VPWR _15280_/X sky130_fd_sc_hd__o21a_4
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12492_ _12503_/A _12492_/B _12491_/Y VGND VGND VPWR VPWR _12492_/X sky130_fd_sc_hd__and3_4
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24478_ _24496_/CLK _24478_/D HRESETn VGND VGND VPWR VPWR _24478_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ _14231_/A VGND VGND VPWR VPWR _14231_/Y sky130_fd_sc_hd__inv_2
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23429_ _23478_/CLK _23429_/D VGND VGND VPWR VPWR _20270_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22445__A2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14162_ _14099_/A _14098_/X _14099_/A _14098_/X VGND VGND VPWR VPWR _14162_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21653__B1 _17722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25263__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13113_ _13113_/A VGND VGND VPWR VPWR _13114_/B sky130_fd_sc_hd__inv_2
X_14093_ _23996_/Q _14078_/A _14073_/X _14023_/A _14076_/A VGND VGND VPWR VPWR _25213_/D
+ sky130_fd_sc_hd__a32o_4
X_18970_ _18969_/Y _14665_/X _17421_/X _14665_/X VGND VGND VPWR VPWR _18970_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22777__A2_N _22773_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_63_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13044_ _12990_/C _13052_/B VGND VGND VPWR VPWR _13045_/B sky130_fd_sc_hd__or2_4
X_17921_ _17921_/A VGND VGND VPWR VPWR _17921_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18787__A _18792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17852_ _17854_/B VGND VGND VPWR VPWR _17853_/B sky130_fd_sc_hd__inv_2
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16803_ _14930_/Y _16797_/X HWDATA[29] _16802_/X VGND VGND VPWR VPWR _16803_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17783_ _17837_/A _17762_/X VGND VGND VPWR VPWR _17786_/B sky130_fd_sc_hd__or2_4
X_14995_ _15166_/B _24461_/Q _14994_/A _24461_/Q VGND VGND VPWR VPWR _14996_/D sky130_fd_sc_hd__a2bb2o_4
X_19522_ _19520_/Y _19516_/X _11939_/X _19521_/X VGND VGND VPWR VPWR _23698_/D sky130_fd_sc_hd__a2bb2o_4
X_16734_ _16739_/A VGND VGND VPWR VPWR _16734_/X sky130_fd_sc_hd__buf_2
X_13946_ _13905_/C _24950_/Q _13945_/X _13946_/D VGND VGND VPWR VPWR _13947_/B sky130_fd_sc_hd__or4_4
XFILLER_130_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22381__B2 _22380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19453_ _19451_/Y _19447_/X _19407_/X _19452_/X VGND VGND VPWR VPWR _23722_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21941__A _17717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16665_ _16662_/Y _16658_/X _16306_/X _16664_/X VGND VGND VPWR VPWR _24489_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19827__A2_N _19824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24145__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13877_ _13871_/X _13876_/X _14268_/A _13867_/X VGND VGND VPWR VPWR _25234_/D sky130_fd_sc_hd__o22a_4
XFILLER_35_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18404_ _18404_/A _18399_/X _18404_/C _18403_/X VGND VGND VPWR VPWR _18404_/X sky130_fd_sc_hd__or4_4
X_15616_ _24888_/Q VGND VGND VPWR VPWR _15616_/Y sky130_fd_sc_hd__inv_2
X_12828_ _25358_/Q VGND VGND VPWR VPWR _12845_/A sky130_fd_sc_hd__inv_2
X_19384_ _19384_/A VGND VGND VPWR VPWR _19384_/X sky130_fd_sc_hd__buf_2
X_16596_ _16594_/Y _16595_/X _16242_/X _16595_/X VGND VGND VPWR VPWR _16596_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18335_ _18334_/X VGND VGND VPWR VPWR _18335_/X sky130_fd_sc_hd__buf_2
X_15547_ _22873_/B VGND VGND VPWR VPWR _15728_/A sky130_fd_sc_hd__buf_2
XANTENNA__12156__A1_N _12092_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12759_ _23181_/A VGND VGND VPWR VPWR _12759_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18266_ _18265_/Y _18262_/Y _16852_/X _18262_/Y VGND VGND VPWR VPWR _18266_/X sky130_fd_sc_hd__a2bb2o_4
X_15478_ _14868_/Y _15476_/X _15477_/X _15476_/X VGND VGND VPWR VPWR _24940_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17217_ _16308_/Y _23008_/A _24609_/Q _17350_/C VGND VGND VPWR VPWR _17224_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14429_ _14428_/Y _14426_/X _14239_/X _14426_/X VGND VGND VPWR VPWR _25126_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15571__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18197_ _18010_/A _23741_/Q VGND VGND VPWR VPWR _18198_/C sky130_fd_sc_hd__or2_4
XANTENNA__19837__B1 _19794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17148_ _17148_/A _17146_/Y _17160_/C VGND VGND VPWR VPWR _17148_/X sky130_fd_sc_hd__and3_4
X_17079_ _16976_/Y _17086_/B VGND VGND VPWR VPWR _17079_/X sky130_fd_sc_hd__or2_4
XFILLER_131_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14721__C _21781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20090_ _20088_/Y _20086_/X _20089_/X _20086_/X VGND VGND VPWR VPWR _20090_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24986__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18697__A _18743_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24915__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22800_ _16823_/A _21067_/A _22797_/X _22799_/X VGND VGND VPWR VPWR _22801_/C sky130_fd_sc_hd__a211o_4
XANTENNA__13634__A _13634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_20_0_HCLK clkbuf_8_21_0_HCLK/A VGND VGND VPWR VPWR _24109_/CLK sky130_fd_sc_hd__clkbuf_1
X_23780_ _23660_/CLK _23780_/D VGND VGND VPWR VPWR _13158_/B sky130_fd_sc_hd__dfxtp_4
X_20992_ _20992_/A _20992_/B VGND VGND VPWR VPWR _20992_/X sky130_fd_sc_hd__and2_4
XANTENNA__17379__A1 _17244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_83_0_HCLK clkbuf_8_83_0_HCLK/A VGND VGND VPWR VPWR _24070_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21851__A _21019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22731_ _22510_/A _22728_/X _22413_/X _22730_/X VGND VGND VPWR VPWR _22731_/X sky130_fd_sc_hd__o22a_4
XFILLER_80_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15929__A2 _15795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22666__B _15854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25450_ _25368_/CLK _12396_/Y HRESETn VGND VGND VPWR VPWR _12266_/A sky130_fd_sc_hd__dfrtp_4
X_22662_ _22659_/X _22662_/B _22661_/X _22658_/A VGND VGND VPWR VPWR _22662_/X sky130_fd_sc_hd__and4_4
XFILLER_111_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24401_ _24998_/CLK _16856_/X HRESETn VGND VGND VPWR VPWR _16855_/A sky130_fd_sc_hd__dfrtp_4
X_21613_ _21609_/X _21612_/X _14749_/X VGND VGND VPWR VPWR _21613_/X sky130_fd_sc_hd__o21a_4
X_25381_ _25368_/CLK _25381_/D HRESETn VGND VGND VPWR VPWR _25381_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_2_3_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_6_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22593_ _21700_/X _22592_/X _21296_/X _24714_/Q _21299_/X VGND VGND VPWR VPWR _22593_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24332_ _24177_/CLK _17375_/Y HRESETn VGND VGND VPWR VPWR _24332_/Q sky130_fd_sc_hd__dfrtp_4
X_21544_ _14393_/Y _14195_/B _14465_/Y _17416_/A VGND VGND VPWR VPWR _21544_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24263_ _24689_/CLK _17824_/X HRESETn VGND VGND VPWR VPWR _24263_/Q sky130_fd_sc_hd__dfrtp_4
X_21475_ _21649_/A _21472_/X _21474_/X VGND VGND VPWR VPWR _21475_/X sky130_fd_sc_hd__and3_4
XANTENNA__22427__A2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23214_ _23034_/X _23213_/X _22466_/X _24870_/Q _23102_/X VGND VGND VPWR VPWR _23214_/X
+ sky130_fd_sc_hd__a32o_4
X_20426_ _20443_/A _20426_/B VGND VGND VPWR VPWR _20428_/C sky130_fd_sc_hd__or2_4
X_24194_ _24186_/CLK _18337_/X HRESETn VGND VGND VPWR VPWR _24194_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13809__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19991__A _19991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23145_ _23034_/X _23144_/X _22968_/X _24868_/Q _23102_/X VGND VGND VPWR VPWR _23145_/X
+ sky130_fd_sc_hd__a32o_4
X_20357_ _20356_/Y _20352_/X _20019_/X _20339_/Y VGND VGND VPWR VPWR _23396_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23076_ _12841_/B _21872_/X _16909_/Y _22821_/X VGND VGND VPWR VPWR _23076_/X sky130_fd_sc_hd__o22a_4
X_20288_ _21786_/B _20283_/X _19988_/X _20283_/X VGND VGND VPWR VPWR _20288_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22027_ _22016_/A _22027_/B VGND VGND VPWR VPWR _22027_/X sky130_fd_sc_hd__or2_4
XFILLER_88_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24656__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16814__B1 _15729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13800_ _16359_/A VGND VGND VPWR VPWR _13800_/X sky130_fd_sc_hd__buf_2
XFILLER_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11992_ _24087_/Q _11992_/B VGND VGND VPWR VPWR _11992_/X sky130_fd_sc_hd__and2_4
X_14780_ _16173_/B VGND VGND VPWR VPWR _14781_/A sky130_fd_sc_hd__inv_2
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18567__B1 _18487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23978_ _23978_/CLK _23978_/D HRESETn VGND VGND VPWR VPWR _17396_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12300__B1 _12299_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21761__A _21616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13731_ _11682_/A _25268_/Q VGND VGND VPWR VPWR _13731_/X sky130_fd_sc_hd__or2_4
XFILLER_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22929_ _22929_/A VGND VGND VPWR VPWR _22929_/X sky130_fd_sc_hd__buf_2
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12585__A2_N _24868_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16450_ _22088_/A VGND VGND VPWR VPWR _16451_/A sky130_fd_sc_hd__buf_2
X_13662_ _24041_/Q _13662_/B VGND VGND VPWR VPWR _13663_/B sky130_fd_sc_hd__or2_4
X_15401_ _15384_/A _15398_/B _15400_/Y VGND VGND VPWR VPWR _24972_/D sky130_fd_sc_hd__and3_4
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ _25398_/Q VGND VGND VPWR VPWR _12712_/A sky130_fd_sc_hd__inv_2
X_13593_ _12049_/A _15782_/B _11714_/Y _13593_/D VGND VGND VPWR VPWR _13593_/X sky130_fd_sc_hd__or4_4
X_16381_ _16381_/A VGND VGND VPWR VPWR _16389_/A sky130_fd_sc_hd__buf_2
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14375__A _11710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18120_ _18005_/A _18118_/X _18120_/C VGND VGND VPWR VPWR _18120_/X sky130_fd_sc_hd__and3_4
XFILLER_101_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12544_ _12534_/X _12537_/X _12540_/X _12543_/X VGND VGND VPWR VPWR _12558_/C sky130_fd_sc_hd__or4_4
X_15332_ _15346_/A _15330_/X _15332_/C VGND VGND VPWR VPWR _24990_/D sky130_fd_sc_hd__and3_4
XANTENNA__25444__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18051_ _17990_/A VGND VGND VPWR VPWR _18187_/A sky130_fd_sc_hd__buf_2
X_12475_ _12475_/A _12475_/B VGND VGND VPWR VPWR _12476_/C sky130_fd_sc_hd__or2_4
X_15263_ _15282_/A _15261_/X _15263_/C VGND VGND VPWR VPWR _15263_/X sky130_fd_sc_hd__and3_4
X_17002_ _16037_/Y _17031_/A _16037_/Y _17031_/A VGND VGND VPWR VPWR _17002_/X sky130_fd_sc_hd__a2bb2o_4
X_14214_ _14214_/A VGND VGND VPWR VPWR _14214_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15194_ _15194_/A _15204_/B VGND VGND VPWR VPWR _15194_/X sky130_fd_sc_hd__or2_4
XANTENNA__18098__A2 _18078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14145_ _14125_/X _14143_/Y _14102_/A _14144_/X VGND VGND VPWR VPWR _25207_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14076_ _14076_/A VGND VGND VPWR VPWR _14076_/X sky130_fd_sc_hd__buf_2
X_18953_ _18951_/Y _18947_/X _17424_/X _18952_/X VGND VGND VPWR VPWR _18953_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21936__A _17706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13027_ _13026_/X VGND VGND VPWR VPWR _25348_/D sky130_fd_sc_hd__inv_2
X_17904_ _17904_/A _17896_/Y VGND VGND VPWR VPWR _17904_/X sky130_fd_sc_hd__or2_4
X_18884_ _18884_/A _18881_/X VGND VGND VPWR VPWR _20562_/A sky130_fd_sc_hd__or2_4
XFILLER_6_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24397__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16805__B1 HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17835_ _17755_/Y _17830_/B _17780_/X _17831_/Y VGND VGND VPWR VPWR _17835_/X sky130_fd_sc_hd__a211o_4
XFILLER_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13454__A _13454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17766_ _17766_/A VGND VGND VPWR VPWR _17768_/B sky130_fd_sc_hd__inv_2
X_14978_ _15166_/C _16799_/A _15166_/C _16799_/A VGND VGND VPWR VPWR _14978_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19505_ _19504_/Y _19500_/X _11948_/X _19500_/X VGND VGND VPWR VPWR _23704_/D sky130_fd_sc_hd__a2bb2o_4
X_16717_ _14470_/A VGND VGND VPWR VPWR _16717_/X sky130_fd_sc_hd__buf_2
X_13929_ _13958_/C VGND VGND VPWR VPWR _13930_/D sky130_fd_sc_hd__buf_2
X_17697_ _17688_/X _17696_/X _17681_/X VGND VGND VPWR VPWR _24279_/D sky130_fd_sc_hd__and3_4
X_19436_ _19435_/Y _19431_/X _19389_/X _19431_/X VGND VGND VPWR VPWR _23728_/D sky130_fd_sc_hd__a2bb2o_4
X_16648_ _16648_/A VGND VGND VPWR VPWR _16648_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22106__A1 _12278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22106__B2 _22821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19367_ _19366_/Y _19361_/X _19232_/X _19361_/X VGND VGND VPWR VPWR _23752_/D sky130_fd_sc_hd__a2bb2o_4
X_16579_ _24519_/Q VGND VGND VPWR VPWR _16579_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23961__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18318_ _18311_/Y _18318_/B _18315_/X _18317_/X VGND VGND VPWR VPWR _18319_/C sky130_fd_sc_hd__or4_4
XANTENNA__21865__B1 _24846_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19298_ _19297_/Y _19295_/X _19206_/X _19295_/X VGND VGND VPWR VPWR _19298_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22933__C _22926_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25114__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18249_ _18249_/A VGND VGND VPWR VPWR _18249_/X sky130_fd_sc_hd__buf_2
XANTENNA__23067__C1 _23066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21260_ _17700_/C VGND VGND VPWR VPWR _21260_/X sky130_fd_sc_hd__buf_2
X_20211_ _20210_/X VGND VGND VPWR VPWR _20211_/Y sky130_fd_sc_hd__inv_2
X_21191_ _21191_/A _21191_/B _21191_/C VGND VGND VPWR VPWR _21191_/X sky130_fd_sc_hd__and3_4
XFILLER_117_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16005__A _24731_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12533__A _12533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15847__A1 _15655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20142_ _23478_/Q VGND VGND VPWR VPWR _20142_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11747__A2_N _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16964__A1_N _16033_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20073_ _20065_/A _18325_/X _20072_/X _23503_/Q _20065_/Y VGND VGND VPWR VPWR _23503_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21565__B _12054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24950_ _24950_/CLK _15455_/X HRESETn VGND VGND VPWR VPWR _24950_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19261__A1_N _21225_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23901_ _24209_/CLK _18943_/X VGND VGND VPWR VPWR _23901_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24067__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24881_ _24883_/CLK _24881_/D HRESETn VGND VGND VPWR VPWR _21280_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23832_ _23832_/CLK _19142_/X VGND VGND VPWR VPWR _18122_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23763_ _23828_/CLK _19337_/X VGND VGND VPWR VPWR _18002_/B sky130_fd_sc_hd__dfxtp_4
X_20975_ _20974_/A _20974_/B _24110_/Q _20974_/X VGND VGND VPWR VPWR _20975_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24500__CLK _23498_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25502_ _25497_/CLK _11907_/X HRESETn VGND VGND VPWR VPWR _11871_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_54_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22714_ _22714_/A VGND VGND VPWR VPWR _22714_/X sky130_fd_sc_hd__buf_2
X_23694_ _23711_/CLK _19531_/X VGND VGND VPWR VPWR _23694_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25433_ _25433_/CLK _25433_/D HRESETn VGND VGND VPWR VPWR _12462_/A sky130_fd_sc_hd__dfrtp_4
X_22645_ _15709_/A _22644_/X _22130_/C _16042_/A _22915_/A VGND VGND VPWR VPWR _22645_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14195__A _14195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20659__A1 _14226_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25364_ _25356_/CLK _25364_/D HRESETn VGND VGND VPWR VPWR _12954_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24650__CLK _24581_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22576_ _22576_/A _22726_/B VGND VGND VPWR VPWR _22576_/X sky130_fd_sc_hd__and2_4
X_21527_ _16640_/A _21526_/X _21427_/X _24809_/Q _21323_/X VGND VGND VPWR VPWR _21528_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_103_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23301__A _24766_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24315_ _24883_/CLK _17433_/X HRESETn VGND VGND VPWR VPWR _24315_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25295_ _25478_/CLK _25295_/D HRESETn VGND VGND VPWR VPWR _13514_/A sky130_fd_sc_hd__dfrtp_4
X_12260_ _12260_/A VGND VGND VPWR VPWR _12433_/A sky130_fd_sc_hd__inv_2
X_24246_ _24248_/CLK _24246_/D HRESETn VGND VGND VPWR VPWR _16926_/A sky130_fd_sc_hd__dfrtp_4
X_21458_ _21458_/A VGND VGND VPWR VPWR _21459_/A sky130_fd_sc_hd__buf_2
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17288__B1 _17236_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20409_ _23374_/Q VGND VGND VPWR VPWR _20409_/Y sky130_fd_sc_hd__inv_2
X_12191_ _12191_/A VGND VGND VPWR VPWR _12290_/A sky130_fd_sc_hd__inv_2
XFILLER_135_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24177_ _24177_/CLK _24177_/D HRESETn VGND VGND VPWR VPWR _21091_/A sky130_fd_sc_hd__dfrtp_4
X_21389_ _21371_/A _20163_/Y VGND VGND VPWR VPWR _21389_/X sky130_fd_sc_hd__or2_4
XANTENNA__12443__A _12440_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24837__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15838__A1 _15824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23128_ _23128_/A _23128_/B VGND VGND VPWR VPWR _23128_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__13849__B1 _13810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15950_ _12207_/Y _15945_/X _15949_/X _15945_/X VGND VGND VPWR VPWR _24759_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23059_ _24557_/Q _22879_/X _22798_/X VGND VGND VPWR VPWR _23059_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24490__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14901_ _25021_/Q VGND VGND VPWR VPWR _15071_/A sky130_fd_sc_hd__inv_2
X_15881_ _12822_/Y _15879_/X _11781_/X _15879_/X VGND VGND VPWR VPWR _15881_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17620_ _17617_/A _17616_/B _17619_/X VGND VGND VPWR VPWR _17620_/X sky130_fd_sc_hd__and3_4
XANTENNA__13274__A _13450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14832_ _14803_/C _14817_/X _14819_/A _14819_/B VGND VGND VPWR VPWR _14832_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15192__C _15171_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14274__B1 _14239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22587__A _24783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11810__A1_N _11807_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21491__A _21491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17551_ _17532_/X _17551_/B _17551_/C _17550_/X VGND VGND VPWR VPWR _17551_/X sky130_fd_sc_hd__or4_4
X_14763_ _13739_/B _14772_/A _14762_/X VGND VGND VPWR VPWR _14763_/X sky130_fd_sc_hd__or3_4
X_11975_ _11647_/X _11970_/C _11974_/X VGND VGND VPWR VPWR _11975_/X sky130_fd_sc_hd__or3_4
XANTENNA__22887__A2 _22523_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16502_ _16501_/Y _16499_/X _16228_/X _16499_/X VGND VGND VPWR VPWR _16502_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13714_ _13714_/A VGND VGND VPWR VPWR _13714_/X sky130_fd_sc_hd__buf_2
X_17482_ _17477_/A VGND VGND VPWR VPWR _17482_/X sky130_fd_sc_hd__buf_2
XFILLER_32_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14694_ _13755_/A _13751_/A _13758_/B VGND VGND VPWR VPWR _14694_/X sky130_fd_sc_hd__a21o_4
X_19221_ _19221_/A VGND VGND VPWR VPWR _19221_/Y sky130_fd_sc_hd__inv_2
X_16433_ _16433_/A VGND VGND VPWR VPWR _16433_/X sky130_fd_sc_hd__buf_2
X_13645_ _25285_/Q _13524_/X _13640_/X VGND VGND VPWR VPWR _13673_/A sky130_fd_sc_hd__a21o_4
XANTENNA__22639__A2 _22821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19152_ _19152_/A _14671_/X _25061_/Q _19152_/D VGND VGND VPWR VPWR _19153_/A sky130_fd_sc_hd__or4_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16364_ _16363_/Y _16282_/A _16266_/X _16282_/A VGND VGND VPWR VPWR _16364_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _13576_/A VGND VGND VPWR VPWR _13576_/Y sky130_fd_sc_hd__inv_2
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _18066_/A _23768_/Q VGND VGND VPWR VPWR _18103_/X sky130_fd_sc_hd__or2_4
X_15315_ _15315_/A VGND VGND VPWR VPWR _15318_/A sky130_fd_sc_hd__buf_2
X_12527_ _12527_/A VGND VGND VPWR VPWR _12527_/Y sky130_fd_sc_hd__inv_2
X_19083_ _19083_/A VGND VGND VPWR VPWR _22361_/B sky130_fd_sc_hd__inv_2
X_16295_ _16295_/A VGND VGND VPWR VPWR _16295_/Y sky130_fd_sc_hd__inv_2
X_18034_ _18168_/A _18034_/B VGND VGND VPWR VPWR _18035_/C sky130_fd_sc_hd__or2_4
X_15246_ _15246_/A VGND VGND VPWR VPWR _15282_/A sky130_fd_sc_hd__buf_2
X_12458_ _12457_/X VGND VGND VPWR VPWR _25434_/D sky130_fd_sc_hd__inv_2
XFILLER_126_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21075__A1 _12983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13449__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12389_ _12389_/A _12389_/B _12389_/C VGND VGND VPWR VPWR _12389_/X sky130_fd_sc_hd__and3_4
X_15177_ _15166_/B _15165_/X VGND VGND VPWR VPWR _15180_/B sky130_fd_sc_hd__or2_4
XANTENNA__24578__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12760__B1 _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14128_ _25131_/Q VGND VGND VPWR VPWR _14128_/Y sky130_fd_sc_hd__inv_2
X_19985_ _11937_/A VGND VGND VPWR VPWR _19985_/X sky130_fd_sc_hd__buf_2
XANTENNA__24507__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19136__A _18996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14059_ _14084_/A VGND VGND VPWR VPWR _14076_/A sky130_fd_sc_hd__buf_2
X_18936_ _13379_/B VGND VGND VPWR VPWR _18936_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18867_ _18866_/X VGND VGND VPWR VPWR _18867_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17818_ _17758_/A _17758_/B _17758_/D _17818_/D VGND VGND VPWR VPWR _17824_/B sky130_fd_sc_hd__or4_4
X_18798_ _18792_/A _18796_/A VGND VGND VPWR VPWR _18798_/X sky130_fd_sc_hd__or2_4
XANTENNA__14265__B1 _13840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17749_ _17748_/Y _16920_/Y _16927_/A VGND VGND VPWR VPWR _17750_/D sky130_fd_sc_hd__or3_4
XFILLER_36_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16495__A _24551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20760_ _20743_/X _20759_/X _24898_/Q _20747_/X VGND VGND VPWR VPWR _20760_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25366__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17002__A1_N _16037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19419_ _19419_/A VGND VGND VPWR VPWR _19419_/Y sky130_fd_sc_hd__inv_2
X_20691_ _20690_/Y _13123_/X _13126_/B VGND VGND VPWR VPWR _20691_/X sky130_fd_sc_hd__o21a_4
XFILLER_50_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_157_0_HCLK clkbuf_7_78_0_HCLK/X VGND VGND VPWR VPWR _24682_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_51_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22430_ _12204_/Y _22407_/B _22266_/X _12318_/Y _21529_/X VGND VGND VPWR VPWR _22430_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__21838__B1 _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23121__A _22786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22361_ _22055_/X _22361_/B VGND VGND VPWR VPWR _22362_/C sky130_fd_sc_hd__or2_4
X_24100_ _23933_/CLK _20965_/X HRESETn VGND VGND VPWR VPWR _24100_/Q sky130_fd_sc_hd__dfrtp_4
X_21312_ _21019_/A VGND VGND VPWR VPWR _21312_/X sky130_fd_sc_hd__buf_2
X_25080_ _25081_/CLK _25080_/D HRESETn VGND VGND VPWR VPWR _14570_/A sky130_fd_sc_hd__dfrtp_4
X_22292_ _23281_/A _22283_/Y _22287_/X _22132_/A _22291_/X VGND VGND VPWR VPWR _22293_/D
+ sky130_fd_sc_hd__o32a_4
XANTENNA__16190__B1 _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23055__A2 _22988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24031_ _24033_/CLK _20827_/Y HRESETn VGND VGND VPWR VPWR _13651_/A sky130_fd_sc_hd__dfrtp_4
X_21243_ _21237_/X _21242_/X _14676_/X VGND VGND VPWR VPWR _21243_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24930__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21174_ _21185_/A _21174_/B VGND VGND VPWR VPWR _21174_/X sky130_fd_sc_hd__or2_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24248__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20125_ _20125_/A VGND VGND VPWR VPWR _22370_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_5_22_0_HCLK_A clkbuf_5_22_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22566__A1 _16898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20056_ _20056_/A VGND VGND VPWR VPWR _20056_/Y sky130_fd_sc_hd__inv_2
X_24933_ _24673_/CLK _15496_/X HRESETn VGND VGND VPWR VPWR _12049_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_86_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24864_ _24847_/CLK _15731_/X HRESETn VGND VGND VPWR VPWR _24864_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23815_ _23832_/CLK _23815_/D VGND VGND VPWR VPWR _19187_/A sky130_fd_sc_hd__dfxtp_4
X_24795_ _24832_/CLK _24795_/D HRESETn VGND VGND VPWR VPWR _24795_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11777_/A VGND VGND VPWR VPWR _11760_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_53_0_HCLK clkbuf_7_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20958_ _12017_/X _20958_/B VGND VGND VPWR VPWR _24090_/D sky130_fd_sc_hd__and2_4
XFILLER_41_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23746_ _23446_/CLK _23746_/D VGND VGND VPWR VPWR _18026_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25036__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _25277_/Q VGND VGND VPWR VPWR _13689_/A sky130_fd_sc_hd__inv_2
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _20889_/A _20889_/B VGND VGND VPWR VPWR _20889_/X sky130_fd_sc_hd__or2_4
X_23677_ _23396_/CLK _23677_/D VGND VGND VPWR VPWR _23677_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ _13177_/Y _13422_/X _13429_/X VGND VGND VPWR VPWR _13430_/X sky130_fd_sc_hd__and3_4
XANTENNA__16226__A1_N _16223_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25416_ _25411_/CLK _12641_/Y HRESETn VGND VGND VPWR VPWR _12606_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22628_ _24611_/Q _22592_/B VGND VGND VPWR VPWR _22628_/X sky130_fd_sc_hd__or2_4
XANTENNA__19498__B2 _19495_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17948__B _19309_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _13453_/A _13361_/B _13361_/C VGND VGND VPWR VPWR _13365_/B sky130_fd_sc_hd__and3_4
XANTENNA__23031__A _24758_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22559_ _22559_/A _22747_/B VGND VGND VPWR VPWR _22559_/X sky130_fd_sc_hd__and2_4
X_25347_ _23370_/CLK _13033_/X HRESETn VGND VGND VPWR VPWR _12299_/A sky130_fd_sc_hd__dfrtp_4
X_15100_ _24971_/Q _24575_/Q _15299_/B _15099_/Y VGND VGND VPWR VPWR _15100_/X sky130_fd_sc_hd__o22a_4
X_12312_ _12311_/Y _24807_/Q _12311_/Y _24807_/Q VGND VGND VPWR VPWR _12312_/X sky130_fd_sc_hd__a2bb2o_4
X_13292_ _13168_/A _13290_/X _13291_/X VGND VGND VPWR VPWR _13292_/X sky130_fd_sc_hd__and3_4
X_16080_ _11739_/A _15655_/A _15927_/X _24701_/Q _16079_/X VGND VGND VPWR VPWR _16080_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_10_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25278_ _25279_/CLK _13711_/X HRESETn VGND VGND VPWR VPWR _25278_/Q sky130_fd_sc_hd__dfrtp_4
X_12243_ _12430_/A _24748_/Q _12430_/A _24748_/Q VGND VGND VPWR VPWR _12243_/X sky130_fd_sc_hd__a2bb2o_4
X_15031_ _25005_/Q VGND VGND VPWR VPWR _15251_/C sky130_fd_sc_hd__inv_2
X_24229_ _23818_/CLK _24229_/D HRESETn VGND VGND VPWR VPWR _24229_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24671__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21486__A _21455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12174_ SSn_S3 _12173_/Y _11862_/X _12173_/Y VGND VGND VPWR VPWR _25453_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24600__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19770_ _13458_/B VGND VGND VPWR VPWR _19770_/Y sky130_fd_sc_hd__inv_2
X_16982_ _24732_/Q _16981_/A _16001_/Y _16981_/Y VGND VGND VPWR VPWR _16989_/A sky130_fd_sc_hd__o22a_4
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18721_ _18738_/A _18721_/B _18721_/C VGND VGND VPWR VPWR _24140_/D sky130_fd_sc_hd__and3_4
XFILLER_7_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15933_ _15933_/A VGND VGND VPWR VPWR _15933_/X sky130_fd_sc_hd__buf_2
XANTENNA__18795__A _18792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17433__B1 _16852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18652_ _18646_/X _18652_/B _18652_/C _18651_/X VGND VGND VPWR VPWR _18667_/B sky130_fd_sc_hd__or4_4
X_15864_ _15864_/A VGND VGND VPWR VPWR _15864_/X sky130_fd_sc_hd__buf_2
XFILLER_76_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14247__B1 _20490_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17603_ _17603_/A VGND VGND VPWR VPWR _24306_/D sky130_fd_sc_hd__inv_2
XFILLER_92_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14815_ _25035_/Q _14814_/X _14815_/C VGND VGND VPWR VPWR _14816_/B sky130_fd_sc_hd__or3_4
XFILLER_36_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18583_ _18475_/B _18559_/X _18581_/B _18498_/X VGND VGND VPWR VPWR _18583_/X sky130_fd_sc_hd__a211o_4
X_15795_ _15795_/A VGND VGND VPWR VPWR _15795_/X sky130_fd_sc_hd__buf_2
XANTENNA__19186__B1 _19117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25119__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17534_ _11770_/Y _24301_/Q _11770_/Y _24301_/Q VGND VGND VPWR VPWR _17537_/B sky130_fd_sc_hd__a2bb2o_4
X_14746_ _14746_/A _14746_/B VGND VGND VPWR VPWR _14746_/X sky130_fd_sc_hd__or2_4
X_11958_ _11957_/Y VGND VGND VPWR VPWR _11958_/X sky130_fd_sc_hd__buf_2
XANTENNA__17736__A1 _17700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18933__B1 _16782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17465_ _24195_/Q VGND VGND VPWR VPWR _17465_/X sky130_fd_sc_hd__buf_2
X_14677_ _14676_/X VGND VGND VPWR VPWR _14677_/X sky130_fd_sc_hd__buf_2
XFILLER_60_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11889_ _11894_/B _11887_/X VGND VGND VPWR VPWR _11889_/Y sky130_fd_sc_hd__nor2_4
X_19204_ _19202_/Y _19198_/X _19136_/X _19203_/X VGND VGND VPWR VPWR _19204_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16416_ _24582_/Q VGND VGND VPWR VPWR _16416_/Y sky130_fd_sc_hd__inv_2
X_13628_ _25061_/Q VGND VGND VPWR VPWR _19014_/A sky130_fd_sc_hd__buf_2
X_17396_ _17396_/A _17396_/B VGND VGND VPWR VPWR _20650_/B sky130_fd_sc_hd__or2_4
XFILLER_38_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19135_ _23834_/Q VGND VGND VPWR VPWR _19135_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16347_ _22402_/A VGND VGND VPWR VPWR _16347_/Y sky130_fd_sc_hd__inv_2
X_13559_ _13559_/A VGND VGND VPWR VPWR _13559_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24759__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19066_ _19065_/Y _19063_/X _18993_/X _19063_/X VGND VGND VPWR VPWR _23859_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16278_ _24630_/Q VGND VGND VPWR VPWR _16278_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18017_ _18017_/A _18017_/B _18016_/X VGND VGND VPWR VPWR _18017_/X sky130_fd_sc_hd__or3_4
X_15229_ _15219_/C _15211_/B _15199_/X _15227_/B VGND VGND VPWR VPWR _15230_/A sky130_fd_sc_hd__a211o_4
XFILLER_114_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19110__B1 _18993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24341__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19968_ _19968_/A VGND VGND VPWR VPWR _19968_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18919_ _19841_/A VGND VGND VPWR VPWR _18919_/X sky130_fd_sc_hd__buf_2
XFILLER_79_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19899_ _23568_/Q VGND VGND VPWR VPWR _21803_/B sky130_fd_sc_hd__inv_2
XFILLER_80_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22939__B _21048_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21930_ _21945_/A _19938_/Y VGND VGND VPWR VPWR _21930_/X sky130_fd_sc_hd__or2_4
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21861_ _23085_/A _21861_/B _21861_/C VGND VGND VPWR VPWR _21861_/X sky130_fd_sc_hd__and3_4
XFILLER_94_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19177__B1 _19155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20812_ _20812_/A VGND VGND VPWR VPWR _20812_/Y sky130_fd_sc_hd__inv_2
X_23600_ _23683_/CLK _19813_/X VGND VGND VPWR VPWR _13363_/B sky130_fd_sc_hd__dfxtp_4
X_21792_ _21456_/A _21792_/B VGND VGND VPWR VPWR _21792_/X sky130_fd_sc_hd__or2_4
X_24580_ _24572_/CLK _16422_/X HRESETn VGND VGND VPWR VPWR _16421_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_36_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20743_ _20770_/A VGND VGND VPWR VPWR _20743_/X sky130_fd_sc_hd__buf_2
XANTENNA__15738__B1 _11791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23531_ _23394_/CLK _23531_/D VGND VGND VPWR VPWR _20004_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23462_ _24089_/CLK _20185_/X VGND VGND VPWR VPWR _23462_/Q sky130_fd_sc_hd__dfxtp_4
X_20674_ _20674_/A VGND VGND VPWR VPWR _20674_/Y sky130_fd_sc_hd__inv_2
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15753__A3 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22413_ _21017_/B VGND VGND VPWR VPWR _22413_/X sky130_fd_sc_hd__buf_2
X_25201_ _25199_/CLK _25201_/D HRESETn VGND VGND VPWR VPWR _14099_/A sky130_fd_sc_hd__dfrtp_4
X_23393_ _23682_/CLK _23393_/D VGND VGND VPWR VPWR _23393_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12972__B1 _12866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22344_ _22025_/A _22342_/X _22343_/X VGND VGND VPWR VPWR _22344_/X sky130_fd_sc_hd__and3_4
XFILLER_52_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25132_ _25093_/CLK _25132_/D HRESETn VGND VGND VPWR VPWR _25132_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__24429__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25063_ _23828_/CLK _25063_/D HRESETn VGND VGND VPWR VPWR _14645_/A sky130_fd_sc_hd__dfrtp_4
X_22275_ _21064_/X _22269_/X _22270_/X _22274_/X VGND VGND VPWR VPWR _22276_/B sky130_fd_sc_hd__a22oi_4
XANTENNA__15910__B1 _24772_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24014_ _24868_/CLK _24014_/D HRESETn VGND VGND VPWR VPWR _13119_/A sky130_fd_sc_hd__dfrtp_4
X_21226_ _21247_/A _21226_/B _21225_/X VGND VGND VPWR VPWR _21226_/X sky130_fd_sc_hd__and3_4
XFILLER_104_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21157_ _15671_/A _21157_/B _21157_/C VGND VGND VPWR VPWR _21157_/X sky130_fd_sc_hd__and3_4
XANTENNA__24011__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20108_ _23491_/Q VGND VGND VPWR VPWR _22209_/B sky130_fd_sc_hd__inv_2
X_21088_ _24632_/Q _15655_/A _21087_/X _21031_/X VGND VGND VPWR VPWR _21089_/A sky130_fd_sc_hd__a211o_4
XFILLER_8_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12440__B _12286_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12930_ _12930_/A VGND VGND VPWR VPWR _12930_/Y sky130_fd_sc_hd__inv_2
X_20039_ _20038_/Y _20036_/X _19995_/X _20036_/X VGND VGND VPWR VPWR _20039_/X sky130_fd_sc_hd__a2bb2o_4
X_24916_ _25255_/CLK _15536_/X HRESETn VGND VGND VPWR VPWR _12057_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_74_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12861_ _12881_/A _12861_/B _12861_/C VGND VGND VPWR VPWR _25386_/D sky130_fd_sc_hd__and3_4
XANTENNA__15977__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24847_ _24847_/CLK _24847_/D HRESETn VGND VGND VPWR VPWR _24847_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19168__B1 _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14600_ _14596_/B _14598_/Y _14599_/X _14590_/X _25076_/Q VGND VGND VPWR VPWR _14600_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_27_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11812_ HWDATA[12] VGND VGND VPWR VPWR _11812_/X sky130_fd_sc_hd__buf_2
XANTENNA__17024__A _17023_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15580_ _15580_/A VGND VGND VPWR VPWR _15588_/A sky130_fd_sc_hd__buf_2
X_12792_ _12792_/A VGND VGND VPWR VPWR _12792_/Y sky130_fd_sc_hd__inv_2
XPHY_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24778_ _24813_/CLK _15903_/X HRESETn VGND VGND VPWR VPWR _24778_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17718__B2 _21465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14521_/X _14530_/X _25102_/Q _14517_/A VGND VGND VPWR VPWR _25090_/D sky130_fd_sc_hd__o22a_4
XPHY_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ HWDATA[31] VGND VGND VPWR VPWR _11743_/X sky130_fd_sc_hd__buf_2
XPHY_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ _23718_/CLK _23729_/D VGND VGND VPWR VPWR _18071_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17250_/A VGND VGND VPWR VPWR _17252_/A sky130_fd_sc_hd__inv_2
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14461_/Y _14459_/X _14391_/X _14459_/X VGND VGND VPWR VPWR _14462_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11673_/Y _24227_/Q _11673_/Y _24227_/Q VGND VGND VPWR VPWR _11675_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_140_0_HCLK clkbuf_7_70_0_HCLK/X VGND VGND VPWR VPWR _25316_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15744__A3 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ _16199_/Y _16200_/X _11761_/X _16200_/X VGND VGND VPWR VPWR _16201_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _13413_/A _13411_/X _13412_/X VGND VGND VPWR VPWR _13414_/C sky130_fd_sc_hd__and3_4
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17181_ _17173_/X _17176_/X _17179_/X _17181_/D VGND VGND VPWR VPWR _17202_/B sky130_fd_sc_hd__or4_4
X_14393_ _14393_/A VGND VGND VPWR VPWR _14393_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24852__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19340__B1 _19294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16132_ _16130_/Y _16126_/X _11804_/X _16131_/X VGND VGND VPWR VPWR _16132_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11800__A _11800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13344_ _13269_/A _23374_/Q VGND VGND VPWR VPWR _13344_/X sky130_fd_sc_hd__or2_4
X_16063_ _24708_/Q VGND VGND VPWR VPWR _16063_/Y sky130_fd_sc_hd__inv_2
X_13275_ _13314_/A _13271_/X _13275_/C VGND VGND VPWR VPWR _13276_/C sky130_fd_sc_hd__or3_4
XANTENNA__15901__B1 _15758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15014_ _25004_/Q _15013_/A _15262_/A _15013_/Y VGND VGND VPWR VPWR _15014_/X sky130_fd_sc_hd__o22a_4
X_12226_ _12215_/X _12218_/X _12222_/X _12226_/D VGND VGND VPWR VPWR _12227_/D sky130_fd_sc_hd__or4_4
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12157_ _12157_/A _12157_/B _12154_/X _12156_/X VGND VGND VPWR VPWR _12157_/X sky130_fd_sc_hd__or4_4
X_19822_ _13736_/X _13762_/X _19822_/C VGND VGND VPWR VPWR _19823_/A sky130_fd_sc_hd__or3_4
XFILLER_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21944__A _21944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12088_ _12088_/A VGND VGND VPWR VPWR _12088_/Y sky130_fd_sc_hd__inv_2
X_16965_ _24370_/Q VGND VGND VPWR VPWR _17041_/D sky130_fd_sc_hd__inv_2
X_19753_ _19749_/Y _19752_/X _19664_/X _19752_/X VGND VGND VPWR VPWR _23620_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15916_ _15685_/X _13588_/X _15677_/A _13590_/A VGND VGND VPWR VPWR _15916_/X sky130_fd_sc_hd__a211o_4
X_18704_ _18704_/A _18703_/X VGND VGND VPWR VPWR _18704_/X sky130_fd_sc_hd__or2_4
XANTENNA__15942__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19684_ _19683_/X VGND VGND VPWR VPWR _19697_/A sky130_fd_sc_hd__inv_2
XFILLER_65_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16896_ _16124_/Y _24261_/Q _16124_/Y _24261_/Q VGND VGND VPWR VPWR _16896_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18635_ _18635_/A _18635_/B _18632_/X _18634_/X VGND VGND VPWR VPWR _18636_/D sky130_fd_sc_hd__or4_4
XFILLER_77_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15847_ _15655_/X _15765_/X _15845_/X _12604_/A _15846_/X VGND VGND VPWR VPWR _24805_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15968__B1 _24751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18566_ _18566_/A _18572_/B VGND VGND VPWR VPWR _18566_/X sky130_fd_sc_hd__or2_4
X_15778_ _15552_/Y _15655_/X _15774_/X _20674_/A _15777_/X VGND VGND VPWR VPWR _15778_/X
+ sky130_fd_sc_hd__a32o_4
X_17517_ _17517_/A VGND VGND VPWR VPWR _17517_/Y sky130_fd_sc_hd__inv_2
X_14729_ _22038_/A _14740_/B VGND VGND VPWR VPWR _14729_/Y sky130_fd_sc_hd__nand2_4
X_18497_ _18457_/Y _18479_/X _18503_/A _18496_/X VGND VGND VPWR VPWR _18497_/X sky130_fd_sc_hd__or4_4
XFILLER_71_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17448_ _11710_/A _17447_/X VGND VGND VPWR VPWR _17448_/X sky130_fd_sc_hd__or2_4
XANTENNA__23258__A2 _21533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17379_ _17244_/Y _17381_/B _17378_/Y VGND VGND VPWR VPWR _17379_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24593__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19118_ _19116_/Y _19112_/X _19117_/X _19112_/X VGND VGND VPWR VPWR _19118_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11710__A _11710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20390_ _20383_/X _20379_/X _18254_/X _23383_/Q _20381_/X VGND VGND VPWR VPWR _23383_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16145__B1 _16143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24522__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19049_ _19049_/A VGND VGND VPWR VPWR _19049_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22060_ _22055_/X _22060_/B VGND VGND VPWR VPWR _22060_/X sky130_fd_sc_hd__or2_4
XFILLER_114_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21011_ _21410_/A VGND VGND VPWR VPWR _22764_/A sky130_fd_sc_hd__buf_2
XFILLER_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21441__A1 _16927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21441__B2 _22429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15852__A _15852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25381__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22962_ _22962_/A VGND VGND VPWR VPWR _23114_/A sky130_fd_sc_hd__buf_2
XANTENNA__22941__A1 _24723_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24701_ _24840_/CLK _16080_/X HRESETn VGND VGND VPWR VPWR _24701_/Q sky130_fd_sc_hd__dfrtp_4
X_21913_ _17717_/A _19502_/Y VGND VGND VPWR VPWR _21916_/B sky130_fd_sc_hd__or2_4
XANTENNA__12293__A2_N _24818_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25310__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22893_ _22759_/X _22892_/X _22854_/X _24826_/Q _22761_/X VGND VGND VPWR VPWR _22894_/B
+ sky130_fd_sc_hd__a32o_4
X_24632_ _24893_/CLK _16274_/X HRESETn VGND VGND VPWR VPWR _24632_/Q sky130_fd_sc_hd__dfrtp_4
X_21844_ _20496_/D _21843_/X _14461_/Y _17416_/A VGND VGND VPWR VPWR _21845_/D sky130_fd_sc_hd__o22a_4
XFILLER_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15974__A3 _11818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21775_ _21771_/X _21774_/X _14749_/X VGND VGND VPWR VPWR _21775_/X sky130_fd_sc_hd__o21a_4
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24563_ _24557_/CLK _16468_/X HRESETn VGND VGND VPWR VPWR _24563_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16683__A _16664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20726_ _20725_/X VGND VGND VPWR VPWR _20726_/X sky130_fd_sc_hd__buf_2
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23514_ _23562_/CLK _23514_/D VGND VGND VPWR VPWR _23514_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24494_ _24492_/CLK _24494_/D HRESETn VGND VGND VPWR VPWR _24494_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15726__A3 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_213_0_HCLK clkbuf_8_213_0_HCLK/A VGND VGND VPWR VPWR _24984_/CLK sky130_fd_sc_hd__clkbuf_1
X_20657_ _20657_/A _20657_/B _20656_/X VGND VGND VPWR VPWR _23980_/D sky130_fd_sc_hd__and3_4
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23445_ _23798_/CLK _20229_/X VGND VGND VPWR VPWR _23445_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16136__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23376_ _24187_/CLK _23376_/D VGND VGND VPWR VPWR _23376_/Q sky130_fd_sc_hd__dfxtp_4
X_20588_ _20587_/X VGND VGND VPWR VPWR _23943_/D sky130_fd_sc_hd__inv_2
XANTENNA__24263__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25115_ _25101_/CLK _14457_/X HRESETn VGND VGND VPWR VPWR _20529_/A sky130_fd_sc_hd__dfrtp_4
X_22327_ _21912_/X _22325_/X _22326_/X VGND VGND VPWR VPWR _22327_/X sky130_fd_sc_hd__and3_4
X_13060_ _13049_/A _13060_/B _13059_/Y VGND VGND VPWR VPWR _25340_/D sky130_fd_sc_hd__and3_4
XFILLER_30_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22258_ _23386_/Q _21995_/Y _22506_/B _22257_/X VGND VGND VPWR VPWR _22259_/A sky130_fd_sc_hd__a211o_4
X_25046_ _23516_/CLK _25046_/D HRESETn VGND VGND VPWR VPWR _25046_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22224__A3 _22219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12011_ _25300_/Q _12010_/Y _25300_/Q _12010_/Y VGND VGND VPWR VPWR _12012_/D sky130_fd_sc_hd__a2bb2o_4
X_21209_ _21209_/A VGND VGND VPWR VPWR _21209_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17019__A _17346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22189_ _22200_/A _22189_/B VGND VGND VPWR VPWR _22189_/X sky130_fd_sc_hd__or2_4
XANTENNA__25469__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21764__A _21616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19474__A2_N _19471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16750_ _15025_/Y _16749_/X _16401_/X _16749_/X VGND VGND VPWR VPWR _24454_/D sky130_fd_sc_hd__a2bb2o_4
X_13962_ _13968_/A _13954_/X _13961_/X VGND VGND VPWR VPWR _13962_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_47_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21735__A2 _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15701_ _15642_/A _15701_/B VGND VGND VPWR VPWR _15702_/A sky130_fd_sc_hd__or2_4
XFILLER_58_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12913_ _12850_/C _12912_/X _12866_/X VGND VGND VPWR VPWR _12913_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__25051__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16681_ _16680_/Y _16676_/X _16325_/X _16676_/X VGND VGND VPWR VPWR _16681_/X sky130_fd_sc_hd__a2bb2o_4
X_13893_ _13927_/A _13893_/B _13953_/A _13947_/A VGND VGND VPWR VPWR _13894_/A sky130_fd_sc_hd__or4_4
XFILLER_47_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18420_ _18420_/A VGND VGND VPWR VPWR _18420_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15632_ _15561_/X VGND VGND VPWR VPWR _15632_/X sky130_fd_sc_hd__buf_2
X_12844_ _25356_/Q VGND VGND VPWR VPWR _12976_/A sky130_fd_sc_hd__inv_2
XFILLER_62_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18792__B _18792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18351_ _18350_/Y _17477_/Y _24187_/Q _17482_/X VGND VGND VPWR VPWR _18365_/B sky130_fd_sc_hd__o22a_4
X_15563_ _15563_/A VGND VGND VPWR VPWR _15563_/X sky130_fd_sc_hd__buf_2
X_12775_ _24779_/Q VGND VGND VPWR VPWR _12775_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_23_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17266_/A _17293_/B _17302_/C VGND VGND VPWR VPWR _24351_/D sky130_fd_sc_hd__and3_4
X_14514_ _20441_/B _14511_/X _14512_/Y _14513_/X VGND VGND VPWR VPWR _14514_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12814__A2_N _24787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _24919_/Q _11726_/B VGND VGND VPWR VPWR _13777_/A sky130_fd_sc_hd__or2_4
X_18282_ _17708_/Y _19492_/B _17709_/Y VGND VGND VPWR VPWR _20276_/C sky130_fd_sc_hd__or3_4
XPHY_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15490_/X VGND VGND VPWR VPWR _15494_/X sky130_fd_sc_hd__buf_2
XPHY_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17233_ _17344_/A VGND VGND VPWR VPWR _17266_/A sky130_fd_sc_hd__buf_2
X_14445_ _14444_/Y _14442_/X _14391_/X _14442_/X VGND VGND VPWR VPWR _14445_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _25279_/Q VGND VGND VPWR VPWR _13691_/A sky130_fd_sc_hd__inv_2
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15002__A _15002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17164_ _17043_/Y _17065_/X _17067_/X _17162_/B VGND VGND VPWR VPWR _17164_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16127__B1 _11796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21939__A _21454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _15991_/A _15991_/B _15991_/C _16369_/D VGND VGND VPWR VPWR _14377_/B sky130_fd_sc_hd__or4_4
XFILLER_70_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12829__A2_N _24775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16115_ _16115_/A VGND VGND VPWR VPWR _16115_/Y sky130_fd_sc_hd__inv_2
X_13327_ _13233_/A VGND VGND VPWR VPWR _13428_/A sky130_fd_sc_hd__buf_2
XANTENNA__17875__B1 _17790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17095_ _16967_/A _17095_/B VGND VGND VPWR VPWR _17095_/X sky130_fd_sc_hd__or2_4
XFILLER_127_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16046_ _24714_/Q VGND VGND VPWR VPWR _16046_/Y sky130_fd_sc_hd__inv_2
X_13258_ _13195_/X VGND VGND VPWR VPWR _13258_/X sky130_fd_sc_hd__buf_2
XFILLER_108_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23986__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12209_ _25427_/Q VGND VGND VPWR VPWR _12209_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13457__A _13457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22620__B1 _22527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13189_ _18344_/A _23908_/Q VGND VGND VPWR VPWR _13189_/X sky130_fd_sc_hd__or2_4
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21974__A2 _20329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19805_ _13253_/B VGND VGND VPWR VPWR _19805_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20949__A1_N _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25139__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17997_ _18080_/A _19020_/A VGND VGND VPWR VPWR _18000_/B sky130_fd_sc_hd__or2_4
X_16948_ _16939_/Y VGND VGND VPWR VPWR _16948_/X sky130_fd_sc_hd__buf_2
X_19736_ _19734_/Y _19730_/X _19645_/X _19735_/X VGND VGND VPWR VPWR _23626_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_105_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_211_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16879_ _16879_/A VGND VGND VPWR VPWR _16879_/Y sky130_fd_sc_hd__inv_2
X_19667_ _19666_/Y _19663_/X _19642_/X _19663_/X VGND VGND VPWR VPWR _19667_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18618_ _24520_/Q _24131_/Q _16577_/Y _18758_/A VGND VGND VPWR VPWR _18625_/A sky130_fd_sc_hd__o22a_4
XFILLER_20_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19598_ _19598_/A VGND VGND VPWR VPWR _19598_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22936__C _23005_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18549_ _18521_/A VGND VGND VPWR VPWR _18555_/A sky130_fd_sc_hd__buf_2
XFILLER_127_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24774__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22151__A2 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14950__A2_N _24415_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21560_ _21559_/X VGND VGND VPWR VPWR _21560_/X sky130_fd_sc_hd__buf_2
XANTENNA__24703__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20511_ _20455_/B _20510_/X _20495_/X VGND VGND VPWR VPWR _20513_/C sky130_fd_sc_hd__o21a_4
X_21491_ _21491_/A _21482_/X _21491_/C VGND VGND VPWR VPWR _21491_/X sky130_fd_sc_hd__or3_4
XFILLER_14_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22952__B _22952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23230_ _20799_/Y _22988_/X _20939_/A _22790_/X VGND VGND VPWR VPWR _23230_/X sky130_fd_sc_hd__o22a_4
X_20442_ _20454_/C VGND VGND VPWR VPWR _20443_/D sky130_fd_sc_hd__inv_2
XFILLER_105_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23161_ _23119_/X _23159_/X _23121_/X _23160_/X VGND VGND VPWR VPWR _23162_/B sky130_fd_sc_hd__o22a_4
X_20373_ _20360_/Y VGND VGND VPWR VPWR _20373_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_43_0_HCLK clkbuf_8_43_0_HCLK/A VGND VGND VPWR VPWR _23869_/CLK sky130_fd_sc_hd__clkbuf_1
X_22112_ _15467_/Y _21352_/X _14228_/Y _14221_/A VGND VGND VPWR VPWR _22112_/X sky130_fd_sc_hd__o22a_4
X_23092_ _23091_/X VGND VGND VPWR VPWR _23092_/Y sky130_fd_sc_hd__inv_2
X_22043_ _22040_/Y _22041_/X _21963_/X _22042_/X VGND VGND VPWR VPWR _22044_/B sky130_fd_sc_hd__a211o_4
XFILLER_86_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24943__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23167__A1 _24560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23994_ _23995_/CLK _20513_/X HRESETn VGND VGND VPWR VPWR _23994_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13814__B _15851_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22945_ _20905_/Y _22824_/X _20767_/A _22280_/A VGND VGND VPWR VPWR _22945_/X sky130_fd_sc_hd__o22a_4
XFILLER_60_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14198__A _14807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19791__B1 _19790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13533__C _15652_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22876_ _20757_/Y _21106_/X _20896_/Y _21211_/X VGND VGND VPWR VPWR _22877_/B sky130_fd_sc_hd__o22a_4
XANTENNA__15947__A3 HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24615_ _24889_/CLK _16326_/X HRESETn VGND VGND VPWR VPWR _24615_/Q sky130_fd_sc_hd__dfrtp_4
X_21827_ _22929_/A VGND VGND VPWR VPWR _22677_/B sky130_fd_sc_hd__buf_2
XANTENNA__22678__B1 _21211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _12560_/A VGND VGND VPWR VPWR _12704_/A sky130_fd_sc_hd__inv_2
XANTENNA__16357__B1 _16355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12091__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24546_ _24465_/CLK _16509_/X HRESETn VGND VGND VPWR VPWR _16508_/A sky130_fd_sc_hd__dfrtp_4
X_21758_ _21754_/X _21757_/X _14749_/X VGND VGND VPWR VPWR _21758_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24444__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20709_ _13129_/A _13129_/B _20708_/Y VGND VGND VPWR VPWR _20709_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_32_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12269_/Y _12491_/B VGND VGND VPWR VPWR _12491_/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24477_ _24041_/CLK _24477_/D HRESETn VGND VGND VPWR VPWR _24477_/Q sky130_fd_sc_hd__dfrtp_4
X_21689_ _21682_/Y _21688_/Y _22035_/A VGND VGND VPWR VPWR _21689_/X sky130_fd_sc_hd__o21a_4
XFILLER_71_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14230_ _14228_/Y _14224_/X _13840_/X _14229_/X VGND VGND VPWR VPWR _14230_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16109__B1 _11771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23428_ _24070_/CLK _20274_/X VGND VGND VPWR VPWR _23428_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22445__A3 _16728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20663__A _20663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14161_ _14146_/X _14160_/Y _25122_/Q _14111_/X VGND VGND VPWR VPWR _25202_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17857__B1 _17790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23359_ _21002_/X VGND VGND VPWR VPWR IRQ[5] sky130_fd_sc_hd__buf_2
X_13112_ _13107_/X _13112_/B _13115_/C VGND VGND VPWR VPWR _25324_/D sky130_fd_sc_hd__and3_4
X_14092_ _14023_/A _20459_/B _14069_/X _14003_/C _14076_/A VGND VGND VPWR VPWR _25214_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_79_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13277__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13043_ _13043_/A _13043_/B VGND VGND VPWR VPWR _13052_/B sky130_fd_sc_hd__or2_4
X_17920_ _17920_/A _17920_/B _17920_/C VGND VGND VPWR VPWR _17921_/A sky130_fd_sc_hd__or3_4
XANTENNA__17972__A _13610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25029_ _25029_/CLK _14879_/Y HRESETn VGND VGND VPWR VPWR _14798_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__12181__A _22267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18787__B _18792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17851_ _16918_/Y _17846_/X _16898_/X _17850_/X VGND VGND VPWR VPWR _17854_/B sky130_fd_sc_hd__or4_4
XANTENNA__25232__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16802_ _16807_/A VGND VGND VPWR VPWR _16802_/X sky130_fd_sc_hd__buf_2
XFILLER_38_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17782_ _17781_/X VGND VGND VPWR VPWR _17782_/Y sky130_fd_sc_hd__inv_2
X_14994_ _14994_/A VGND VGND VPWR VPWR _15166_/B sky130_fd_sc_hd__buf_2
XFILLER_59_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22102__B _21105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16733_ _16733_/A VGND VGND VPWR VPWR _16739_/A sky130_fd_sc_hd__buf_2
X_19521_ _19528_/A VGND VGND VPWR VPWR _19521_/X sky130_fd_sc_hd__buf_2
X_13945_ _13945_/A _13905_/A _13901_/X VGND VGND VPWR VPWR _13945_/X sky130_fd_sc_hd__or3_4
XFILLER_47_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22381__A2 _22352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19452_ _19446_/Y VGND VGND VPWR VPWR _19452_/X sky130_fd_sc_hd__buf_2
XFILLER_75_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16664_ _16664_/A VGND VGND VPWR VPWR _16664_/X sky130_fd_sc_hd__buf_2
XFILLER_62_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13876_ _21716_/A _13860_/X _25233_/Q _13855_/X VGND VGND VPWR VPWR _13876_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16596__B1 _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15615_ _22513_/A _15612_/X _11825_/X _15612_/X VGND VGND VPWR VPWR _15615_/X sky130_fd_sc_hd__a2bb2o_4
X_18403_ _16268_/Y _24145_/Q _16268_/Y _24145_/Q VGND VGND VPWR VPWR _18403_/X sky130_fd_sc_hd__a2bb2o_4
X_12827_ _12817_/X _12827_/B _12823_/X _12826_/X VGND VGND VPWR VPWR _12827_/X sky130_fd_sc_hd__or4_4
X_19383_ _18026_/B VGND VGND VPWR VPWR _19383_/Y sky130_fd_sc_hd__inv_2
X_16595_ _16583_/A VGND VGND VPWR VPWR _16595_/X sky130_fd_sc_hd__buf_2
X_18334_ _17467_/Y _17449_/X VGND VGND VPWR VPWR _18334_/X sky130_fd_sc_hd__or2_4
XFILLER_128_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15546_ _22915_/A VGND VGND VPWR VPWR _22873_/B sky130_fd_sc_hd__buf_2
XANTENNA__12082__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12758_ _22967_/A VGND VGND VPWR VPWR _12758_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16348__B1 _16057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24185__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14555__B _14555_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11709_ _11707_/Y _11709_/B VGND VGND VPWR VPWR _11710_/A sky130_fd_sc_hd__or2_4
X_18265_ _18265_/A VGND VGND VPWR VPWR _18265_/Y sky130_fd_sc_hd__inv_2
X_15477_ _15986_/A VGND VGND VPWR VPWR _15477_/X sky130_fd_sc_hd__buf_2
XANTENNA__24114__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12689_ _12686_/A _12689_/B _12689_/C VGND VGND VPWR VPWR _12689_/X sky130_fd_sc_hd__and3_4
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17216_ _17212_/X _17213_/X _17214_/X _17215_/X VGND VGND VPWR VPWR _17216_/X sky130_fd_sc_hd__or4_4
XFILLER_129_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14428_ _25126_/Q VGND VGND VPWR VPWR _14428_/Y sky130_fd_sc_hd__inv_2
X_18196_ _18196_/A _18196_/B VGND VGND VPWR VPWR _18198_/B sky130_fd_sc_hd__or2_4
X_17147_ _17020_/X VGND VGND VPWR VPWR _17160_/C sky130_fd_sc_hd__buf_2
XANTENNA__21644__A1 _18272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14359_ _25147_/Q _14351_/X _25146_/Q _14356_/X VGND VGND VPWR VPWR _14359_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22841__B1 _12341_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_2_0_HCLK clkbuf_8_3_0_HCLK/A VGND VGND VPWR VPWR _23434_/CLK sky130_fd_sc_hd__clkbuf_1
X_17078_ _17048_/A _17077_/X VGND VGND VPWR VPWR _17086_/B sky130_fd_sc_hd__or2_4
XFILLER_104_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16029_ _16029_/A VGND VGND VPWR VPWR _16029_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20080__B1 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19719_ _19719_/A VGND VGND VPWR VPWR _19719_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20991_ _24324_/Q _20990_/B _24323_/Q _20990_/X VGND VGND VPWR VPWR _20991_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24955__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22730_ _17252_/A _22419_/X _22729_/Y VGND VGND VPWR VPWR _22730_/X sky130_fd_sc_hd__o21a_4
XFILLER_4_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15929__A3 _15927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22661_ _12430_/A _21524_/X _17759_/A _22425_/X VGND VGND VPWR VPWR _22661_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23321__B2 _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24400_ _24398_/CLK _16860_/X HRESETn VGND VGND VPWR VPWR _20079_/A sky130_fd_sc_hd__dfrtp_4
X_21612_ _21612_/A _21610_/X _21611_/X VGND VGND VPWR VPWR _21612_/X sky130_fd_sc_hd__and3_4
XANTENNA__17122__A _17036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25380_ _25368_/CLK _25380_/D HRESETn VGND VGND VPWR VPWR _12749_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_21_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22592_ _16336_/A _22592_/B VGND VGND VPWR VPWR _22592_/X sky130_fd_sc_hd__or2_4
XFILLER_21_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24331_ _24330_/CLK _17379_/X HRESETn VGND VGND VPWR VPWR _24331_/Q sky130_fd_sc_hd__dfrtp_4
X_21543_ _14425_/Y _14223_/A _14169_/Y _15462_/A VGND VGND VPWR VPWR _21543_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21474_ _21670_/A _20313_/Y VGND VGND VPWR VPWR _21474_/X sky130_fd_sc_hd__or2_4
X_24262_ _24689_/CLK _17827_/X HRESETn VGND VGND VPWR VPWR _17826_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22427__A3 _22422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20425_ _20445_/B _20424_/Y VGND VGND VPWR VPWR _20425_/X sky130_fd_sc_hd__and2_4
XANTENNA__12376__B2 _24811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23213_ _23213_/A _23101_/B VGND VGND VPWR VPWR _23213_/X sky130_fd_sc_hd__or2_4
XANTENNA__14481__A _14481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24193_ _24197_/CLK _18341_/X HRESETn VGND VGND VPWR VPWR _13177_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_134_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20356_ _23396_/Q VGND VGND VPWR VPWR _20356_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23144_ _24798_/Q _23101_/B VGND VGND VPWR VPWR _23144_/X sky130_fd_sc_hd__or2_4
XFILLER_66_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23075_ _22646_/A _23075_/B _23074_/X VGND VGND VPWR VPWR _23075_/X sky130_fd_sc_hd__and3_4
X_20287_ _23423_/Q VGND VGND VPWR VPWR _21786_/B sky130_fd_sc_hd__inv_2
XANTENNA__16502__A1_N _16501_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22026_ _22022_/X _22025_/X _21679_/X VGND VGND VPWR VPWR _22026_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_102_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23018__B _22832_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16517__A1_N _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11991_ _11991_/A _11991_/B VGND VGND VPWR VPWR _11992_/B sky130_fd_sc_hd__and2_4
XANTENNA__24696__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23977_ _23978_/CLK _23977_/D HRESETn VGND VGND VPWR VPWR _20642_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19764__B1 _19740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13730_ _13683_/B _13729_/Y _13680_/X _13714_/A _25270_/Q VGND VGND VPWR VPWR _25270_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_84_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22928_ _15096_/A _23171_/B VGND VGND VPWR VPWR _22932_/B sky130_fd_sc_hd__or2_4
XFILLER_95_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16578__B1 _16408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24625__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13661_ _24040_/Q _13661_/B VGND VGND VPWR VPWR _13662_/B sky130_fd_sc_hd__or2_4
X_22859_ _22897_/A _22859_/B VGND VGND VPWR VPWR _22868_/C sky130_fd_sc_hd__and2_4
X_15400_ _15299_/A _15400_/B VGND VGND VPWR VPWR _15400_/Y sky130_fd_sc_hd__nand2_4
X_12612_ _12708_/A _12707_/A _12706_/A _12595_/Y VGND VGND VPWR VPWR _12612_/X sky130_fd_sc_hd__or4_4
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16380_ HWDATA[29] VGND VGND VPWR VPWR _16380_/X sky130_fd_sc_hd__buf_2
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13592_ _14619_/A _13591_/Y VGND VGND VPWR VPWR _13634_/A sky130_fd_sc_hd__or2_4
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15331_ _15331_/A _15329_/A VGND VGND VPWR VPWR _15332_/C sky130_fd_sc_hd__or2_4
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12543_ _25395_/Q _12542_/A _12706_/A _12542_/Y VGND VGND VPWR VPWR _12543_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17967__A _18024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21874__A1 _25424_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24529_ _24553_/CLK _16556_/X HRESETn VGND VGND VPWR VPWR _24529_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22592__B _22592_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24198__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18050_ _18150_/A _23834_/Q VGND VGND VPWR VPWR _18053_/B sky130_fd_sc_hd__or2_4
XFILLER_40_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15262_ _15262_/A _15262_/B VGND VGND VPWR VPWR _15263_/C sky130_fd_sc_hd__or2_4
XFILLER_8_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12474_ _12474_/A _12474_/B VGND VGND VPWR VPWR _12476_/B sky130_fd_sc_hd__or2_4
XANTENNA__16750__B1 _16401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17001_ _16031_/Y _24377_/Q _24724_/Q _17035_/A VGND VGND VPWR VPWR _17001_/X sky130_fd_sc_hd__a2bb2o_4
X_14213_ _14212_/Y _14210_/X _13515_/X _14201_/A VGND VGND VPWR VPWR _14213_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12367__B2 _12366_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15193_ _15193_/A _15193_/B VGND VGND VPWR VPWR _15204_/B sky130_fd_sc_hd__or2_4
XANTENNA__14391__A _16355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25484__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12904__A _12851_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14144_ _14125_/A VGND VGND VPWR VPWR _14144_/X sky130_fd_sc_hd__buf_2
XFILLER_10_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16502__B1 _16228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25413__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18798__A _18792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14075_ _13997_/X _14065_/X _14057_/X _13989_/X _14066_/X VGND VGND VPWR VPWR _25225_/D
+ sky130_fd_sc_hd__a32o_4
X_18952_ _18946_/Y VGND VGND VPWR VPWR _18952_/X sky130_fd_sc_hd__buf_2
X_13026_ _13026_/A _13026_/B _13025_/X VGND VGND VPWR VPWR _13026_/X sky130_fd_sc_hd__or3_4
X_17903_ _17900_/B _17889_/X VGND VGND VPWR VPWR _17905_/A sky130_fd_sc_hd__or2_4
X_18883_ _18882_/Y VGND VGND VPWR VPWR _18883_/X sky130_fd_sc_hd__buf_2
XFILLER_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20062__B1 _19841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17834_ _17834_/A _17832_/X _17834_/C VGND VGND VPWR VPWR _24260_/D sky130_fd_sc_hd__and3_4
XANTENNA__23000__B1 _22997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14977_ _25025_/Q VGND VGND VPWR VPWR _15166_/C sky130_fd_sc_hd__inv_2
X_17765_ _16916_/Y _16948_/X _17765_/C _17765_/D VGND VGND VPWR VPWR _17766_/A sky130_fd_sc_hd__or4_4
X_19504_ _23704_/Q VGND VGND VPWR VPWR _19504_/Y sky130_fd_sc_hd__inv_2
X_13928_ _13946_/D _13909_/X VGND VGND VPWR VPWR _13958_/C sky130_fd_sc_hd__or2_4
X_16716_ _16716_/A VGND VGND VPWR VPWR _16716_/Y sky130_fd_sc_hd__inv_2
X_17696_ _17527_/A _17696_/B VGND VGND VPWR VPWR _17696_/X sky130_fd_sc_hd__or2_4
XANTENNA__24366__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16647_ _23285_/A _16646_/X _16285_/X _16646_/X VGND VGND VPWR VPWR _24496_/D sky130_fd_sc_hd__a2bb2o_4
X_19435_ _18108_/B VGND VGND VPWR VPWR _19435_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13859_ _13851_/A _13857_/X _13852_/X _13858_/Y VGND VGND VPWR VPWR _25240_/D sky130_fd_sc_hd__a211o_4
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22106__A2 _15784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16578_ _16577_/Y _16575_/X _16408_/X _16575_/X VGND VGND VPWR VPWR _16578_/X sky130_fd_sc_hd__a2bb2o_4
X_19366_ _23752_/Q VGND VGND VPWR VPWR _19366_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22783__A _22783_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15529_ _15535_/A VGND VGND VPWR VPWR _15529_/X sky130_fd_sc_hd__buf_2
X_18317_ _18280_/X _18316_/X _18280_/A _18316_/X VGND VGND VPWR VPWR _18317_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17877__A _16927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21865__A1 _24776_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19297_ _13319_/B VGND VGND VPWR VPWR _19297_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21865__B2 _21067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16781__A HWDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18248_ _18235_/X _18237_/X _18247_/X _24220_/Q _18238_/X VGND VGND VPWR VPWR _18248_/X
+ sky130_fd_sc_hd__a32o_4
X_18179_ _18211_/A _19032_/A VGND VGND VPWR VPWR _18181_/B sky130_fd_sc_hd__or2_4
XFILLER_116_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20210_ _25059_/Q _14670_/X _14656_/Y _18987_/D VGND VGND VPWR VPWR _20210_/X sky130_fd_sc_hd__or4_4
X_21190_ _21185_/A _20018_/Y VGND VGND VPWR VPWR _21191_/C sky130_fd_sc_hd__or2_4
XANTENNA__22290__B2 _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18606__A1_N _16581_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20141_ _21629_/B _20140_/X _20096_/X _20140_/X VGND VGND VPWR VPWR _20141_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_117_0_HCLK clkbuf_7_58_0_HCLK/X VGND VGND VPWR VPWR _24555_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18246__B1 _16604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20072_ _11856_/X VGND VGND VPWR VPWR _20072_/X sky130_fd_sc_hd__buf_2
XANTENNA__23119__A _22783_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20053__B1 _19787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12530__B2 _24842_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23900_ _23905_/CLK _23900_/D VGND VGND VPWR VPWR _18944_/A sky130_fd_sc_hd__dfxtp_4
X_24880_ _24893_/CLK _24880_/D HRESETn VGND VGND VPWR VPWR _24880_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16021__A _24724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16272__A2 _15993_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23831_ _25264_/CLK _19145_/X VGND VGND VPWR VPWR _23831_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15860__A _23035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22677__B _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23762_ _23828_/CLK _23762_/D VGND VGND VPWR VPWR _18045_/B sky130_fd_sc_hd__dfxtp_4
X_20974_ _20974_/A _20974_/B VGND VGND VPWR VPWR _20974_/X sky130_fd_sc_hd__and2_4
XFILLER_96_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25501_ _25497_/CLK _11913_/X HRESETn VGND VGND VPWR VPWR _11878_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22396__C _22396_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22713_ _16130_/Y _22426_/X _22712_/X _11802_/Y _22271_/X VGND VGND VPWR VPWR _22713_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__14476__A _14481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24036__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23693_ _23396_/CLK _19533_/X VGND VGND VPWR VPWR _19532_/A sky130_fd_sc_hd__dfxtp_4
X_25432_ _25449_/CLK _25432_/D HRESETn VGND VGND VPWR VPWR _25432_/Q sky130_fd_sc_hd__dfrtp_4
X_22644_ _24612_/Q _22644_/B VGND VGND VPWR VPWR _22644_/X sky130_fd_sc_hd__or2_4
XANTENNA__22648__A3 _22130_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12597__B2 _24845_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25363_ _25356_/CLK _25363_/D HRESETn VGND VGND VPWR VPWR _25363_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22575_ _22575_/A VGND VGND VPWR VPWR _22726_/B sky130_fd_sc_hd__buf_2
X_24314_ _24883_/CLK _17435_/X HRESETn VGND VGND VPWR VPWR _24314_/Q sky130_fd_sc_hd__dfrtp_4
X_21526_ _21526_/A _22879_/A VGND VGND VPWR VPWR _21526_/X sky130_fd_sc_hd__or2_4
XFILLER_21_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16732__B1 _15714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25294_ _25478_/CLK _25294_/D HRESETn VGND VGND VPWR VPWR _25294_/Q sky130_fd_sc_hd__dfrtp_4
X_24245_ _24248_/CLK _24245_/D HRESETn VGND VGND VPWR VPWR _21048_/A sky130_fd_sc_hd__dfrtp_4
X_21457_ _18307_/X VGND VGND VPWR VPWR _21458_/A sky130_fd_sc_hd__buf_2
XFILLER_120_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12190_ _22550_/A VGND VGND VPWR VPWR _12190_/Y sky130_fd_sc_hd__inv_2
X_20408_ _20407_/Y _20405_/X _15766_/X _20405_/X VGND VGND VPWR VPWR _23375_/D sky130_fd_sc_hd__a2bb2o_4
X_21388_ _21388_/A _21388_/B _21387_/X VGND VGND VPWR VPWR _21388_/X sky130_fd_sc_hd__or3_4
XFILLER_107_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24176_ _24171_/CLK _18485_/X HRESETn VGND VGND VPWR VPWR _24176_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_13_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_23127_ _20786_/Y _22988_/X _20925_/Y _22790_/X VGND VGND VPWR VPWR _23128_/B sky130_fd_sc_hd__o22a_4
X_20339_ _20338_/X VGND VGND VPWR VPWR _20339_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_76_0_HCLK clkbuf_6_38_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_76_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22033__A1 _21681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23058_ _16207_/A _23057_/X VGND VGND VPWR VPWR _23058_/X sky130_fd_sc_hd__or2_4
XFILLER_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24877__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14900_ _14900_/A VGND VGND VPWR VPWR _14900_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22584__A2 _22422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22009_ _22009_/A VGND VGND VPWR VPWR _22024_/A sky130_fd_sc_hd__buf_2
XFILLER_62_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15880_ _12758_/Y _15879_/X _11778_/X _15879_/X VGND VGND VPWR VPWR _15880_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18252__A3 _15836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24806__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14831_ _14831_/A VGND VGND VPWR VPWR _23987_/D sky130_fd_sc_hd__buf_2
XFILLER_64_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17550_ _17550_/A _17550_/B _17550_/C _17549_/X VGND VGND VPWR VPWR _17550_/X sky130_fd_sc_hd__or4_4
X_14762_ _25046_/Q _25045_/Q _14762_/C VGND VGND VPWR VPWR _14762_/X sky130_fd_sc_hd__and3_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11974_ _11701_/A _11701_/B _11880_/Y VGND VGND VPWR VPWR _11974_/X sky130_fd_sc_hd__o21a_4
X_16501_ _16501_/A VGND VGND VPWR VPWR _16501_/Y sky130_fd_sc_hd__inv_2
X_13713_ _13713_/A VGND VGND VPWR VPWR _13714_/A sky130_fd_sc_hd__buf_2
X_17481_ _17476_/A _17449_/X _17481_/C VGND VGND VPWR VPWR _17481_/X sky130_fd_sc_hd__and3_4
X_14693_ _14693_/A VGND VGND VPWR VPWR _21612_/A sky130_fd_sc_hd__buf_2
XFILLER_32_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16432_ _15105_/Y _16429_/X _16057_/X _16429_/X VGND VGND VPWR VPWR _16432_/X sky130_fd_sc_hd__a2bb2o_4
X_19220_ _19105_/A _18331_/X _19219_/X VGND VGND VPWR VPWR _19221_/A sky130_fd_sc_hd__or3_4
XANTENNA__11803__A HWDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13644_ _13644_/A VGND VGND VPWR VPWR _13644_/X sky130_fd_sc_hd__buf_2
XANTENNA__24475__CLK _24581_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23297__B1 _22797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12618__B _12565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19151_ _23828_/Q VGND VGND VPWR VPWR _19151_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13785__B1 _13472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16363_ _24600_/Q VGND VGND VPWR VPWR _16363_/Y sky130_fd_sc_hd__inv_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _13575_/A VGND VGND VPWR VPWR _13575_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18102_ _18023_/X _18102_/B _18101_/X VGND VGND VPWR VPWR _18102_/X sky130_fd_sc_hd__and3_4
XFILLER_40_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ _15346_/A _15314_/B _15314_/C VGND VGND VPWR VPWR _15314_/X sky130_fd_sc_hd__and3_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ _12526_/A VGND VGND VPWR VPWR _12526_/Y sky130_fd_sc_hd__inv_2
X_19082_ _19081_/Y _19076_/X _19010_/X _19062_/Y VGND VGND VPWR VPWR _19082_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23049__B1 _12896_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16294_ _16293_/Y _16289_/X _15944_/X _16289_/X VGND VGND VPWR VPWR _16294_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18033_ _17982_/X _18033_/B VGND VGND VPWR VPWR _18033_/X sky130_fd_sc_hd__or2_4
XANTENNA__13537__B1 _13472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15245_ _15245_/A VGND VGND VPWR VPWR _15245_/Y sky130_fd_sc_hd__inv_2
X_12457_ _12238_/X _12430_/X _12402_/X _12454_/B VGND VGND VPWR VPWR _12457_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16106__A _16094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15176_ _15176_/A VGND VGND VPWR VPWR _25025_/D sky130_fd_sc_hd__inv_2
X_12388_ _12179_/Y _12385_/X VGND VGND VPWR VPWR _12389_/C sky130_fd_sc_hd__or2_4
XFILLER_119_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14127_ _14097_/A _14103_/X _14119_/C _14106_/B VGND VGND VPWR VPWR _14127_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19984_ _19984_/A VGND VGND VPWR VPWR _21938_/B sky130_fd_sc_hd__inv_2
XFILLER_114_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14058_ _14056_/A VGND VGND VPWR VPWR _14084_/A sky130_fd_sc_hd__inv_2
X_18935_ _18934_/Y _18930_/X _16787_/X _18930_/X VGND VGND VPWR VPWR _18935_/X sky130_fd_sc_hd__a2bb2o_4
X_13009_ _13001_/X _13017_/D _12374_/Y VGND VGND VPWR VPWR _13009_/X sky130_fd_sc_hd__o21a_4
X_18866_ _18823_/Y _18724_/A _18844_/X _18865_/X VGND VGND VPWR VPWR _18866_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24547__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17817_ _17817_/A VGND VGND VPWR VPWR _17817_/Y sky130_fd_sc_hd__inv_2
X_18797_ _18630_/A _18796_/Y VGND VGND VPWR VPWR _18797_/X sky130_fd_sc_hd__or2_4
XANTENNA__16776__A _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17748_ _24248_/Q VGND VGND VPWR VPWR _17748_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22869__A1_N _12199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21535__B1 _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17679_ _17652_/X _17676_/B _17679_/C VGND VGND VPWR VPWR _17679_/X sky130_fd_sc_hd__and3_4
XFILLER_63_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19418_ _19417_/Y _19415_/X _19349_/X _19415_/X VGND VGND VPWR VPWR _23734_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20690_ _24000_/Q VGND VGND VPWR VPWR _20690_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21838__A1 _24506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19349_ _19055_/X VGND VGND VPWR VPWR _19349_/X sky130_fd_sc_hd__buf_2
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22360_ _14682_/B _19262_/Y VGND VGND VPWR VPWR _22360_/X sky130_fd_sc_hd__or2_4
XANTENNA__25335__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21311_ _15125_/A _22927_/A VGND VGND VPWR VPWR _21320_/B sky130_fd_sc_hd__or2_4
X_22291_ _25361_/Q _22288_/X _22290_/X VGND VGND VPWR VPWR _22291_/X sky130_fd_sc_hd__a21o_4
X_21242_ _21238_/X _21239_/X _21241_/X VGND VGND VPWR VPWR _21242_/X sky130_fd_sc_hd__and3_4
X_24030_ _24035_/CLK _20823_/Y HRESETn VGND VGND VPWR VPWR _24030_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20761__A _20761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21173_ _21173_/A VGND VGND VPWR VPWR _21185_/A sky130_fd_sc_hd__buf_2
XANTENNA__15855__A _15854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20124_ _20122_/Y _20118_/X _20123_/X _20105_/X VGND VGND VPWR VPWR _23485_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24970__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22566__A2 _22425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20055_ _20054_/Y _20050_/X _19790_/X _20050_/X VGND VGND VPWR VPWR _23512_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14889__A1_N _14888_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24932_ _24248_/CLK _15497_/X HRESETn VGND VGND VPWR VPWR _15782_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_24_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24288__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24863_ _24427_/CLK _24863_/D HRESETn VGND VGND VPWR VPWR _12526_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23814_ _23832_/CLK _19192_/X VGND VGND VPWR VPWR _18189_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24498__CLK _23498_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12267__B1 _12266_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24794_ _24792_/CLK _15878_/X HRESETn VGND VGND VPWR VPWR _24794_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _23772_/CLK _23745_/D VGND VGND VPWR VPWR _23745_/Q sky130_fd_sc_hd__dfxtp_4
X_20957_ _11997_/B _20958_/B VGND VGND VPWR VPWR _24089_/D sky130_fd_sc_hd__and2_4
XFILLER_96_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12522__A2_N _24858_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11689_/Y _24213_/Q _11689_/Y _24213_/Q VGND VGND VPWR VPWR _11690_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23676_ _23384_/CLK _19589_/X VGND VGND VPWR VPWR _22385_/A sky130_fd_sc_hd__dfxtp_4
X_20888_ _20889_/A VGND VGND VPWR VPWR _20888_/Y sky130_fd_sc_hd__inv_2
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25415_ _25400_/CLK _12646_/X HRESETn VGND VGND VPWR VPWR _25415_/Q sky130_fd_sc_hd__dfrtp_4
X_22627_ _22476_/X _22626_/X _21285_/A _24819_/Q _22551_/X VGND VGND VPWR VPWR _22627_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13360_ _13392_/A _13360_/B VGND VGND VPWR VPWR _13361_/C sky130_fd_sc_hd__or2_4
XANTENNA__25076__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25346_ _23370_/CLK _13035_/X HRESETn VGND VGND VPWR VPWR _25346_/Q sky130_fd_sc_hd__dfrtp_4
X_22558_ _22544_/X _22556_/X _22125_/X _25517_/Q _22922_/A VGND VGND VPWR VPWR _22558_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16705__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12311_ _25322_/Q VGND VGND VPWR VPWR _12311_/Y sky130_fd_sc_hd__inv_2
X_21509_ _21494_/Y _21506_/Y _22035_/A VGND VGND VPWR VPWR _21509_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25005__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13291_ _13395_/A _19807_/A VGND VGND VPWR VPWR _13291_/X sky130_fd_sc_hd__or2_4
X_25277_ _25279_/CLK _25277_/D HRESETn VGND VGND VPWR VPWR _25277_/Q sky130_fd_sc_hd__dfrtp_4
X_22489_ _22489_/A VGND VGND VPWR VPWR _22489_/X sky130_fd_sc_hd__buf_2
X_15030_ _24450_/Q VGND VGND VPWR VPWR _15030_/Y sky130_fd_sc_hd__inv_2
X_12242_ _12242_/A VGND VGND VPWR VPWR _12430_/A sky130_fd_sc_hd__buf_2
X_24228_ _24346_/CLK _18234_/X HRESETn VGND VGND VPWR VPWR _11664_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12173_ _12173_/A VGND VGND VPWR VPWR _12173_/Y sky130_fd_sc_hd__inv_2
X_24159_ _24159_/CLK _18548_/Y HRESETn VGND VGND VPWR VPWR _24159_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16981_ _16981_/A VGND VGND VPWR VPWR _16981_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20017__B1 _19995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18720_ _18696_/A _18717_/X VGND VGND VPWR VPWR _18721_/C sky130_fd_sc_hd__or2_4
Xclkbuf_8_100_0_HCLK clkbuf_7_50_0_HCLK/X VGND VGND VPWR VPWR _25172_/CLK sky130_fd_sc_hd__clkbuf_1
X_15932_ _15967_/A VGND VGND VPWR VPWR _15933_/A sky130_fd_sc_hd__buf_2
XFILLER_7_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24640__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_163_0_HCLK clkbuf_7_81_0_HCLK/X VGND VGND VPWR VPWR _23580_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_37_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_6_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15863_ _15863_/A VGND VGND VPWR VPWR _15864_/A sky130_fd_sc_hd__buf_2
X_18651_ _16585_/Y _18767_/A _16585_/Y _18767_/A VGND VGND VPWR VPWR _18651_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14814_ _14799_/C _14813_/X _14814_/C VGND VGND VPWR VPWR _14814_/X sky130_fd_sc_hd__or3_4
X_17602_ _17559_/A _17600_/X _17601_/X _17596_/B VGND VGND VPWR VPWR _17603_/A sky130_fd_sc_hd__a211o_4
XFILLER_114_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15794_ _15781_/X _15788_/X _15553_/X _24838_/Q _15793_/X VGND VGND VPWR VPWR _15794_/X
+ sky130_fd_sc_hd__a32o_4
X_18582_ _18562_/B _18582_/B _18582_/C VGND VGND VPWR VPWR _24150_/D sky130_fd_sc_hd__and3_4
XFILLER_33_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14745_ _14744_/X VGND VGND VPWR VPWR _14746_/B sky130_fd_sc_hd__inv_2
X_17533_ _11807_/Y _24291_/Q _11807_/Y _24291_/Q VGND VGND VPWR VPWR _17533_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11957_ _25539_/Q VGND VGND VPWR VPWR _11957_/Y sky130_fd_sc_hd__inv_2
X_17464_ _13174_/X _17453_/B _17456_/Y VGND VGND VPWR VPWR _17472_/B sky130_fd_sc_hd__o21a_4
XANTENNA__19700__A _19055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14676_ _14676_/A VGND VGND VPWR VPWR _14676_/X sky130_fd_sc_hd__buf_2
X_11888_ _11869_/X VGND VGND VPWR VPWR _11894_/B sky130_fd_sc_hd__inv_2
X_16415_ _16412_/Y _16414_/X _16325_/X _16414_/X VGND VGND VPWR VPWR _16415_/X sky130_fd_sc_hd__a2bb2o_4
X_19203_ _19197_/X VGND VGND VPWR VPWR _19203_/X sky130_fd_sc_hd__buf_2
X_13627_ _13609_/X _14792_/A _13623_/Y _13626_/X VGND VGND VPWR VPWR _13627_/X sky130_fd_sc_hd__or4_4
XANTENNA__23222__A _23281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17395_ _20642_/A _20642_/B VGND VGND VPWR VPWR _17396_/B sky130_fd_sc_hd__or2_4
X_16346_ _16345_/Y _16343_/X _16147_/X _16343_/X VGND VGND VPWR VPWR _16346_/X sky130_fd_sc_hd__a2bb2o_4
X_19134_ _19132_/Y _19130_/X _19133_/X _19130_/X VGND VGND VPWR VPWR _23835_/D sky130_fd_sc_hd__a2bb2o_4
X_13558_ _13557_/Y _14559_/A _13557_/Y _14559_/A VGND VGND VPWR VPWR _13558_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12509_ _12509_/A _12509_/B _12509_/C VGND VGND VPWR VPWR _12509_/X sky130_fd_sc_hd__and3_4
X_19065_ _13204_/B VGND VGND VPWR VPWR _19065_/Y sky130_fd_sc_hd__inv_2
X_16277_ _15669_/X _15993_/Y _16270_/X _24631_/Q _16276_/X VGND VGND VPWR VPWR _24631_/D
+ sky130_fd_sc_hd__a32o_4
X_13489_ _13476_/Y VGND VGND VPWR VPWR _13489_/X sky130_fd_sc_hd__buf_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15228_ _15216_/A _15228_/B _15228_/C VGND VGND VPWR VPWR _25012_/D sky130_fd_sc_hd__and3_4
X_18016_ _18057_/A _18013_/X _18015_/X VGND VGND VPWR VPWR _18016_/X sky130_fd_sc_hd__and3_4
XANTENNA__14183__B1 _14182_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24799__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15159_ _15153_/Y VGND VGND VPWR VPWR _15159_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18051__A _17990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24728__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19967_ _19966_/Y _19964_/X _19632_/X _19964_/X VGND VGND VPWR VPWR _19967_/X sky130_fd_sc_hd__a2bb2o_4
X_18918_ _23909_/Q VGND VGND VPWR VPWR _18918_/Y sky130_fd_sc_hd__inv_2
X_19898_ _21937_/B _19895_/X _19622_/X _19895_/X VGND VGND VPWR VPWR _19898_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24381__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22953__C1 _22952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18849_ _18845_/X _18849_/B _18849_/C _18849_/D VGND VGND VPWR VPWR _18849_/X sky130_fd_sc_hd__or4_4
XFILLER_28_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22301__A _23170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24310__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21860_ _24405_/Q _21858_/X _21556_/X _21859_/X VGND VGND VPWR VPWR _21861_/C sky130_fd_sc_hd__a211o_4
X_20811_ _20674_/A _24028_/Q _13137_/X _23318_/A _20725_/X VGND VGND VPWR VPWR _24028_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_93_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21791_ _21787_/X _21790_/X _17722_/X VGND VGND VPWR VPWR _21799_/B sky130_fd_sc_hd__o21a_4
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23530_ _23714_/CLK _23530_/D VGND VGND VPWR VPWR _20006_/A sky130_fd_sc_hd__dfxtp_4
X_20742_ _20721_/X _20741_/X _24894_/Q _20726_/X VGND VGND VPWR VPWR _20742_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25516__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23461_ _24089_/CLK _20187_/X VGND VGND VPWR VPWR _20186_/A sky130_fd_sc_hd__dfxtp_4
X_20673_ _20602_/X _20504_/B VGND VGND VPWR VPWR _20673_/X sky130_fd_sc_hd__and2_4
XFILLER_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23276__A3 _21514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22116__A1_N _14205_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25200_ _25199_/CLK _25200_/D HRESETn VGND VGND VPWR VPWR _14098_/D sky130_fd_sc_hd__dfrtp_4
X_22412_ _22287_/A _22411_/X VGND VGND VPWR VPWR _22412_/X sky130_fd_sc_hd__and2_4
X_23392_ _23714_/CLK _23392_/D VGND VGND VPWR VPWR _20368_/A sky130_fd_sc_hd__dfxtp_4
X_25131_ _25113_/CLK _25131_/D HRESETn VGND VGND VPWR VPWR _25131_/Q sky130_fd_sc_hd__dfstp_4
X_22343_ _22005_/X _19608_/Y VGND VGND VPWR VPWR _22343_/X sky130_fd_sc_hd__or2_4
XANTENNA__21587__A _21408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25062_ _23722_/CLK _14655_/X HRESETn VGND VGND VPWR VPWR _25062_/Q sky130_fd_sc_hd__dfrtp_4
X_22274_ _22271_/X _22273_/X _21290_/C _24709_/Q _21067_/X VGND VGND VPWR VPWR _22274_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_3_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15910__B2 _15864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24013_ _24018_/CLK _24013_/D HRESETn VGND VGND VPWR VPWR _13119_/C sky130_fd_sc_hd__dfrtp_4
X_21225_ _21249_/A _21225_/B VGND VGND VPWR VPWR _21225_/X sky130_fd_sc_hd__or2_4
XANTENNA__24469__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21156_ _16792_/Y _15852_/Y _21314_/A _21155_/X VGND VGND VPWR VPWR _21157_/C sky130_fd_sc_hd__a211o_4
XANTENNA__18860__B1 _21837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25125__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20107_ _22364_/B _20106_/X _20079_/X _20106_/X VGND VGND VPWR VPWR _20107_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25188__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21087_ _21003_/A _21074_/B VGND VGND VPWR VPWR _21087_/X sky130_fd_sc_hd__and2_4
XFILLER_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12440__C _12440_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20038_ _20038_/A VGND VGND VPWR VPWR _20038_/Y sky130_fd_sc_hd__inv_2
X_24915_ _25255_/CLK _15537_/X HRESETn VGND VGND VPWR VPWR _12068_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23307__A _24630_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_236_0_HCLK clkbuf_8_237_0_HCLK/A VGND VGND VPWR VPWR _24813_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_37_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24051__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12860_ _12744_/Y _12858_/A VGND VGND VPWR VPWR _12861_/C sky130_fd_sc_hd__or2_4
XFILLER_46_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24846_ _24842_/CLK _24846_/D HRESETn VGND VGND VPWR VPWR _24846_/Q sky130_fd_sc_hd__dfrtp_4
X_11811_ _25519_/Q VGND VGND VPWR VPWR _11811_/Y sky130_fd_sc_hd__inv_2
X_12791_ _12791_/A _12763_/X _12791_/C _12790_/X VGND VGND VPWR VPWR _12791_/X sky130_fd_sc_hd__or4_4
XPHY_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24777_ _24780_/CLK _24777_/D HRESETn VGND VGND VPWR VPWR _24777_/Q sky130_fd_sc_hd__dfrtp_4
X_21989_ _21989_/A VGND VGND VPWR VPWR _21989_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _21334_/A _14510_/X _21119_/A _14505_/X VGND VGND VPWR VPWR _14530_/X sky130_fd_sc_hd__o22a_4
XPHY_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11741_/X VGND VGND VPWR VPWR _11742_/X sky130_fd_sc_hd__buf_2
XFILLER_15_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23728_ _23718_/CLK _23728_/D VGND VGND VPWR VPWR _18108_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__25257__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _25113_/Q VGND VGND VPWR VPWR _14461_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _13693_/D VGND VGND VPWR VPWR _11673_/Y sky130_fd_sc_hd__inv_2
XPHY_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23659_ _23635_/CLK _23659_/D VGND VGND VPWR VPWR _13242_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _16217_/A VGND VGND VPWR VPWR _16200_/X sky130_fd_sc_hd__buf_2
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _13312_/A _13412_/B VGND VGND VPWR VPWR _13412_/X sky130_fd_sc_hd__or2_4
X_17180_ _16365_/Y _17242_/A _16365_/Y _17242_/A VGND VGND VPWR VPWR _17181_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14392_ _20496_/D _14382_/X _14391_/X _14384_/X VGND VGND VPWR VPWR _14392_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16131_ _16125_/X VGND VGND VPWR VPWR _16131_/X sky130_fd_sc_hd__buf_2
XFILLER_70_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13343_ _13173_/X _13339_/X _13342_/X VGND VGND VPWR VPWR _13343_/X sky130_fd_sc_hd__or3_4
X_25329_ _25351_/CLK _25329_/D HRESETn VGND VGND VPWR VPWR _25329_/Q sky130_fd_sc_hd__dfrtp_4
X_16062_ _16059_/Y _16060_/X _16061_/X _16060_/X VGND VGND VPWR VPWR _16062_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24327__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13274_ _13450_/A _13272_/X _13274_/C VGND VGND VPWR VPWR _13275_/C sky130_fd_sc_hd__and3_4
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24892__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15013_ _15013_/A VGND VGND VPWR VPWR _15013_/Y sky130_fd_sc_hd__inv_2
X_12225_ _25422_/Q _21526_/A _12499_/A _12224_/Y VGND VGND VPWR VPWR _12226_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17103__B1 _17056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20789__B2 _20774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24821__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19821_ _19821_/A VGND VGND VPWR VPWR _22353_/B sky130_fd_sc_hd__inv_2
X_12156_ _12092_/Y _12155_/X _12092_/Y _12155_/X VGND VGND VPWR VPWR _12156_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24139__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12631__B _12631_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_46_0_HCLK clkbuf_6_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_93_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19752_ _19751_/Y VGND VGND VPWR VPWR _19752_/X sky130_fd_sc_hd__buf_2
X_12087_ _12085_/Y _12086_/X _11858_/X _12086_/X VGND VGND VPWR VPWR _25468_/D sky130_fd_sc_hd__a2bb2o_4
X_16964_ _16033_/Y _17030_/A _16033_/Y _17030_/A VGND VGND VPWR VPWR _16964_/X sky130_fd_sc_hd__a2bb2o_4
X_18703_ _18772_/A _18669_/A VGND VGND VPWR VPWR _18703_/X sky130_fd_sc_hd__and2_4
X_15915_ _25289_/Q _15915_/B VGND VGND VPWR VPWR _15915_/X sky130_fd_sc_hd__and2_4
X_19683_ _19683_/A _19683_/B _19683_/C VGND VGND VPWR VPWR _19683_/X sky130_fd_sc_hd__or3_4
X_16895_ _16890_/X _16895_/B _16893_/X _16895_/D VGND VGND VPWR VPWR _16895_/X sky130_fd_sc_hd__or4_4
XANTENNA__22121__A _24777_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20410__B1 _15768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18634_ _16618_/A _18633_/A _16618_/Y _18682_/B VGND VGND VPWR VPWR _18634_/X sky130_fd_sc_hd__o22a_4
X_15846_ _15777_/B _15703_/A VGND VGND VPWR VPWR _15846_/X sky130_fd_sc_hd__or2_4
XFILLER_91_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18565_ _18416_/Y _18574_/B VGND VGND VPWR VPWR _18572_/B sky130_fd_sc_hd__or2_4
X_12989_ _13054_/A _13061_/A _12989_/C VGND VGND VPWR VPWR _12990_/C sky130_fd_sc_hd__or3_4
X_15777_ _15777_/A _15777_/B VGND VGND VPWR VPWR _15777_/X sky130_fd_sc_hd__or2_4
XFILLER_45_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_HCLK clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17516_ _25536_/Q _17515_/A _11748_/Y _17597_/A VGND VGND VPWR VPWR _17516_/X sky130_fd_sc_hd__o22a_4
X_14728_ _14727_/Y _14707_/Y _22036_/A _14707_/A VGND VGND VPWR VPWR _14740_/B sky130_fd_sc_hd__o22a_4
X_18496_ _18496_/A _18772_/A VGND VGND VPWR VPWR _18496_/X sky130_fd_sc_hd__and2_4
XFILLER_127_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14659_ _14659_/A _14659_/B VGND VGND VPWR VPWR _14659_/X sky130_fd_sc_hd__or2_4
X_17447_ _12049_/A _15640_/B _11716_/A _13593_/D VGND VGND VPWR VPWR _17447_/X sky130_fd_sc_hd__or4_4
XANTENNA__18046__A _18046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17378_ _17244_/Y _17381_/B _17271_/X VGND VGND VPWR VPWR _17378_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_53_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19117_ _16786_/X VGND VGND VPWR VPWR _19117_/X sky130_fd_sc_hd__buf_2
XFILLER_9_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16329_ _22703_/A VGND VGND VPWR VPWR _16329_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17342__B1 _17289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24909__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19048_ _19047_/Y _19045_/X _18955_/X _19045_/X VGND VGND VPWR VPWR _23865_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20229__B1 _19771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24562__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21010_ _21009_/X VGND VGND VPWR VPWR _21410_/A sky130_fd_sc_hd__inv_2
XANTENNA__21441__A2 _22821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18842__B1 _16506_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22961_ _22938_/X _22942_/X _22961_/C _22961_/D VGND VGND VPWR VPWR HRDATA[20] sky130_fd_sc_hd__or4_4
XANTENNA__20401__B1 _18247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24700_ _24700_/CLK _24700_/D HRESETn VGND VGND VPWR VPWR _24700_/Q sky130_fd_sc_hd__dfrtp_4
X_21912_ _21194_/A VGND VGND VPWR VPWR _21912_/X sky130_fd_sc_hd__buf_2
XANTENNA__22941__A2 _21021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15481__A1_N _14881_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22892_ _22892_/A _23140_/B VGND VGND VPWR VPWR _22892_/X sky130_fd_sc_hd__or2_4
XFILLER_55_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24631_ _24893_/CLK _24631_/D HRESETn VGND VGND VPWR VPWR _24631_/Q sky130_fd_sc_hd__dfrtp_4
X_21843_ _14192_/X VGND VGND VPWR VPWR _21843_/X sky130_fd_sc_hd__buf_2
XFILLER_83_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12269__A _25426_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_66_0_HCLK clkbuf_8_67_0_HCLK/A VGND VGND VPWR VPWR _25093_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25350__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24562_ _24561_/CLK _24562_/D HRESETn VGND VGND VPWR VPWR _16469_/A sky130_fd_sc_hd__dfrtp_4
X_21774_ _21631_/A _21772_/X _21774_/C VGND VGND VPWR VPWR _21774_/X sky130_fd_sc_hd__and3_4
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23513_ _25264_/CLK _20053_/X VGND VGND VPWR VPWR _23513_/Q sky130_fd_sc_hd__dfxtp_4
X_20725_ _20747_/A VGND VGND VPWR VPWR _20725_/X sky130_fd_sc_hd__buf_2
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24493_ _24413_/CLK _24493_/D HRESETn VGND VGND VPWR VPWR _16653_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23444_ _23660_/CLK _20234_/X VGND VGND VPWR VPWR _13183_/B sky130_fd_sc_hd__dfxtp_4
X_20656_ _23980_/Q _17398_/B _20655_/Y _20604_/Y VGND VGND VPWR VPWR _20656_/X sky130_fd_sc_hd__a211o_4
XFILLER_11_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22457__B2 _22271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23375_ _24187_/CLK _23375_/D VGND VGND VPWR VPWR _23375_/Q sky130_fd_sc_hd__dfxtp_4
X_20587_ _14128_/Y _20556_/A _20546_/X _20586_/Y VGND VGND VPWR VPWR _20587_/X sky130_fd_sc_hd__a211o_4
XFILLER_104_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23947__D sda_i_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25114_ _25113_/CLK _25114_/D HRESETn VGND VGND VPWR VPWR _14458_/A sky130_fd_sc_hd__dfrtp_4
X_22326_ _21458_/A _20275_/Y VGND VGND VPWR VPWR _22326_/X sky130_fd_sc_hd__or2_4
XFILLER_30_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15895__B1 _24783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25045_ _23516_/CLK _25045_/D HRESETn VGND VGND VPWR VPWR _25045_/Q sky130_fd_sc_hd__dfrtp_4
X_22257_ _21978_/B _19585_/A VGND VGND VPWR VPWR _22257_/X sky130_fd_sc_hd__and2_4
XFILLER_105_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12010_ _12010_/A VGND VGND VPWR VPWR _12010_/Y sky130_fd_sc_hd__inv_2
X_21208_ _21127_/X _21138_/X _21208_/C _21207_/X VGND VGND VPWR VPWR _21208_/X sky130_fd_sc_hd__and4_4
X_22188_ _21381_/A VGND VGND VPWR VPWR _22200_/A sky130_fd_sc_hd__buf_2
XFILLER_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24232__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21139_ _14275_/Y _21139_/B VGND VGND VPWR VPWR _21139_/X sky130_fd_sc_hd__or2_4
XFILLER_59_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13961_ _13960_/A _13959_/Y _13960_/Y _13958_/X VGND VGND VPWR VPWR _13961_/X sky130_fd_sc_hd__o22a_4
XFILLER_47_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12912_ _12764_/Y _12850_/B _12753_/X _12903_/X VGND VGND VPWR VPWR _12912_/X sky130_fd_sc_hd__or4_4
X_15700_ _12050_/X _11719_/B _15700_/C _15991_/D VGND VGND VPWR VPWR _15701_/B sky130_fd_sc_hd__or4_4
X_16680_ _24482_/Q VGND VGND VPWR VPWR _16680_/Y sky130_fd_sc_hd__inv_2
X_13892_ _13892_/A VGND VGND VPWR VPWR _13947_/A sky130_fd_sc_hd__buf_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25438__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16072__B1 _15986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12843_ _12843_/A VGND VGND VPWR VPWR _12944_/C sky130_fd_sc_hd__inv_2
X_15631_ _24883_/Q VGND VGND VPWR VPWR _21739_/A sky130_fd_sc_hd__inv_2
X_24829_ _24852_/CLK _15808_/X HRESETn VGND VGND VPWR VPWR _12368_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22145__B1 _25512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12179__A _25451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15562_ _15561_/X VGND VGND VPWR VPWR _15563_/A sky130_fd_sc_hd__buf_2
X_18350_ _24187_/Q VGND VGND VPWR VPWR _18350_/Y sky130_fd_sc_hd__inv_2
X_12774_ _25362_/Q VGND VGND VPWR VPWR _12774_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22696__A1 _24415_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25091__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14513_/A VGND VGND VPWR VPWR _14513_/X sky130_fd_sc_hd__buf_2
X_17301_ _17237_/A _17304_/B VGND VGND VPWR VPWR _17302_/C sky130_fd_sc_hd__or2_4
XFILLER_37_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _13813_/A _11725_/B VGND VGND VPWR VPWR _11733_/A sky130_fd_sc_hd__or2_4
XFILLER_70_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25020__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _15549_/A _15491_/X HADDR[23] _15491_/X VGND VGND VPWR VPWR _15493_/X sky130_fd_sc_hd__a2bb2o_4
X_18281_ _17702_/A VGND VGND VPWR VPWR _19492_/B sky130_fd_sc_hd__buf_2
XANTENNA__14394__A _14394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12907__A _25376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _25121_/Q VGND VGND VPWR VPWR _14444_/Y sky130_fd_sc_hd__inv_2
X_17232_ _17231_/X VGND VGND VPWR VPWR _17344_/A sky130_fd_sc_hd__buf_2
XANTENNA__22448__A1 _16249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _11656_/A VGND VGND VPWR VPWR _11656_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17163_ _17159_/B _17163_/B _17160_/C VGND VGND VPWR VPWR _17163_/X sky130_fd_sc_hd__and3_4
XANTENNA__22999__A2 _22998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14375_ _11710_/A VGND VGND VPWR VPWR _15642_/A sky130_fd_sc_hd__buf_2
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21120__B2 _21355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16114_ _16112_/Y _16113_/X _15955_/X _16113_/X VGND VGND VPWR VPWR _16114_/X sky130_fd_sc_hd__a2bb2o_4
X_13326_ _13453_/A _13324_/X _13325_/X VGND VGND VPWR VPWR _13326_/X sky130_fd_sc_hd__and3_4
X_17094_ _17093_/X VGND VGND VPWR VPWR _17095_/B sky130_fd_sc_hd__inv_2
X_16045_ _16044_/Y _16040_/X _11813_/X _16040_/X VGND VGND VPWR VPWR _16045_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21020__A _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13257_ _13200_/X _13231_/X _13256_/X _25320_/Q _11965_/X VGND VGND VPWR VPWR _13257_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__12353__A2_N _24820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12208_ _12206_/A _12207_/A _12277_/B _12207_/Y VGND VGND VPWR VPWR _12208_/X sky130_fd_sc_hd__o22a_4
X_13188_ _13188_/A _13186_/X _13188_/C VGND VGND VPWR VPWR _13188_/X sky130_fd_sc_hd__and3_4
XFILLER_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19804_ _19801_/Y _19803_/X _18247_/X _19803_/X VGND VGND VPWR VPWR _19804_/X sky130_fd_sc_hd__a2bb2o_4
X_12139_ _12138_/X VGND VGND VPWR VPWR _12139_/Y sky130_fd_sc_hd__inv_2
X_17996_ _17996_/A VGND VGND VPWR VPWR _18080_/A sky130_fd_sc_hd__buf_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19735_ _19729_/Y VGND VGND VPWR VPWR _19735_/X sky130_fd_sc_hd__buf_2
X_16947_ _16090_/Y _24275_/Q _16090_/Y _24275_/Q VGND VGND VPWR VPWR _16947_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23955__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19666_ _23651_/Q VGND VGND VPWR VPWR _19666_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16878_ _20096_/A VGND VGND VPWR VPWR _16879_/A sky130_fd_sc_hd__buf_2
XFILLER_64_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22786__A _22786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18617_ _24131_/Q VGND VGND VPWR VPWR _18758_/A sky130_fd_sc_hd__inv_2
XANTENNA__21690__A _21539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15829_ _15829_/A VGND VGND VPWR VPWR _15829_/X sky130_fd_sc_hd__buf_2
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25108__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19597_ _19597_/A VGND VGND VPWR VPWR _19598_/A sky130_fd_sc_hd__buf_2
XFILLER_92_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15810__B1 _11778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19001__B1 _18955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18548_ _18548_/A VGND VGND VPWR VPWR _18548_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17599__B _17837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18479_ _18458_/Y _18442_/Y _18479_/C _18478_/X VGND VGND VPWR VPWR _18479_/X sky130_fd_sc_hd__or4_4
X_20510_ _20447_/A _20443_/D VGND VGND VPWR VPWR _20510_/X sky130_fd_sc_hd__and2_4
X_21490_ _21485_/X _21489_/X _18299_/X VGND VGND VPWR VPWR _21491_/C sky130_fd_sc_hd__o21a_4
XFILLER_14_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20441_ _20441_/A _20441_/B _20441_/C VGND VGND VPWR VPWR _20454_/C sky130_fd_sc_hd__or3_4
XFILLER_118_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17315__B1 _17279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24743__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23160_ _15572_/Y _23052_/B VGND VGND VPWR VPWR _23160_/X sky130_fd_sc_hd__and2_4
X_20372_ _23390_/Q VGND VGND VPWR VPWR _20372_/Y sky130_fd_sc_hd__inv_2
X_22111_ _22111_/A _22111_/B VGND VGND VPWR VPWR _22111_/X sky130_fd_sc_hd__and2_4
X_23091_ _22753_/X _23089_/X _22684_/X _23090_/X VGND VGND VPWR VPWR _23091_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16024__A _24723_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12552__A _12552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22042_ _14734_/Y _19598_/A VGND VGND VPWR VPWR _22042_/X sky130_fd_sc_hd__and2_4
XANTENNA__15892__A3 _11809_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18815__B1 _18707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21584__B _21019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23993_ _23978_/CLK _20450_/X HRESETn VGND VGND VPWR VPWR _23993_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19240__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22944_ _12433_/A _22820_/X _22943_/X VGND VGND VPWR VPWR _22944_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_112_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25531__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22875_ _23054_/A _22875_/B VGND VGND VPWR VPWR _22875_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15801__B1 _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24614_ _24889_/CLK _16328_/X HRESETn VGND VGND VPWR VPWR _24614_/Q sky130_fd_sc_hd__dfrtp_4
X_21826_ _21826_/A VGND VGND VPWR VPWR _21826_/X sky130_fd_sc_hd__buf_2
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22678__A1 _21106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21105__A _21105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24545_ _24545_/CLK _16512_/X HRESETn VGND VGND VPWR VPWR _16510_/A sky130_fd_sc_hd__dfrtp_4
X_21757_ _21612_/A _21757_/B _21757_/C VGND VGND VPWR VPWR _21757_/X sky130_fd_sc_hd__and3_4
XFILLER_12_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20708_ _20707_/X VGND VGND VPWR VPWR _20708_/Y sky130_fd_sc_hd__inv_2
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12490_ _12209_/Y _12492_/B _12489_/Y VGND VGND VPWR VPWR _12490_/X sky130_fd_sc_hd__o21a_4
X_24476_ _24041_/CLK _24476_/D HRESETn VGND VGND VPWR VPWR _24476_/Q sky130_fd_sc_hd__dfrtp_4
X_21688_ _21687_/X VGND VGND VPWR VPWR _21688_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23320__A _22782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23427_ _23394_/CLK _23427_/D VGND VGND VPWR VPWR _23427_/Q sky130_fd_sc_hd__dfxtp_4
X_20639_ _20642_/B _20638_/Y _20651_/C VGND VGND VPWR VPWR _20639_/X sky130_fd_sc_hd__and3_4
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24484__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18414__A _18414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14160_ _14159_/X VGND VGND VPWR VPWR _14160_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17857__A1 _16898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23358_ _20984_/X VGND VGND VPWR VPWR IRQ[4] sky130_fd_sc_hd__buf_2
XFILLER_4_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24413__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13111_ _13107_/A _13106_/X VGND VGND VPWR VPWR _13112_/B sky130_fd_sc_hd__nand2_4
XFILLER_125_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22309_ _22302_/Y _22309_/B _22309_/C _22308_/Y VGND VGND VPWR VPWR _22309_/X sky130_fd_sc_hd__or4_4
X_14091_ _14063_/X VGND VGND VPWR VPWR _20459_/B sky130_fd_sc_hd__buf_2
Xclkbuf_7_111_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_223_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_23289_ _20807_/Y _22280_/X _20946_/Y _22790_/X VGND VGND VPWR VPWR _23289_/X sky130_fd_sc_hd__o22a_4
X_13042_ _13042_/A VGND VGND VPWR VPWR _13049_/A sky130_fd_sc_hd__buf_2
X_25028_ _23989_/CLK _14883_/Y HRESETn VGND VGND VPWR VPWR _14870_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15773__A HWDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17850_ _16911_/Y _17867_/A _16928_/Y _17850_/D VGND VGND VPWR VPWR _17850_/X sky130_fd_sc_hd__or4_4
XFILLER_105_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18787__C _18608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16801_ _16801_/A VGND VGND VPWR VPWR _16807_/A sky130_fd_sc_hd__buf_2
X_17781_ _16948_/X _17771_/X _17780_/X _17776_/Y VGND VGND VPWR VPWR _17781_/X sky130_fd_sc_hd__a211o_4
X_14993_ _25023_/Q VGND VGND VPWR VPWR _14994_/A sky130_fd_sc_hd__inv_2
XFILLER_120_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19520_ _23698_/Q VGND VGND VPWR VPWR _19520_/Y sky130_fd_sc_hd__inv_2
X_16732_ _15017_/Y _16730_/X _15714_/X _16730_/X VGND VGND VPWR VPWR _16732_/X sky130_fd_sc_hd__a2bb2o_4
X_13944_ _13943_/X VGND VGND VPWR VPWR _13944_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25272__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16045__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19451_ _18036_/B VGND VGND VPWR VPWR _19451_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13875_ _13871_/X _13874_/X _14266_/A _13867_/X VGND VGND VPWR VPWR _13875_/X sky130_fd_sc_hd__o22a_4
X_16663_ _16643_/Y VGND VGND VPWR VPWR _16664_/A sky130_fd_sc_hd__buf_2
XANTENNA__25201__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18402_ _22992_/A _18400_/Y _23200_/A _18503_/A VGND VGND VPWR VPWR _18404_/C sky130_fd_sc_hd__a2bb2o_4
X_12826_ _25377_/Q _12824_/Y _12849_/D _24792_/Q VGND VGND VPWR VPWR _12826_/X sky130_fd_sc_hd__a2bb2o_4
X_15614_ _15614_/A VGND VGND VPWR VPWR _22513_/A sky130_fd_sc_hd__inv_2
X_19382_ _19381_/Y _19379_/X _19291_/X _19379_/X VGND VGND VPWR VPWR _19382_/X sky130_fd_sc_hd__a2bb2o_4
X_16594_ _16594_/A VGND VGND VPWR VPWR _16594_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18333_ _17465_/X VGND VGND VPWR VPWR _18333_/X sky130_fd_sc_hd__buf_2
XANTENNA__21015__A _21015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12757_ _12843_/A _12755_/Y _12854_/A _24798_/Q VGND VGND VPWR VPWR _12757_/X sky130_fd_sc_hd__a2bb2o_4
X_15545_ _15544_/X VGND VGND VPWR VPWR _22915_/A sky130_fd_sc_hd__buf_2
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _24065_/Q VGND VGND VPWR VPWR _11709_/B sky130_fd_sc_hd__inv_2
X_15476_ _15476_/A VGND VGND VPWR VPWR _15476_/X sky130_fd_sc_hd__buf_2
X_18264_ _13795_/D _18253_/X _18254_/X _24211_/Q _18262_/A VGND VGND VPWR VPWR _24211_/D
+ sky130_fd_sc_hd__a32o_4
X_12688_ _25403_/Q _12688_/B VGND VGND VPWR VPWR _12689_/C sky130_fd_sc_hd__or2_4
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ _14425_/Y _14426_/X _14395_/X _14426_/X VGND VGND VPWR VPWR _14427_/X sky130_fd_sc_hd__a2bb2o_4
X_17215_ _16327_/Y _17250_/A _16327_/Y _17250_/A VGND VGND VPWR VPWR _17215_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19298__B1 _19206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18195_ _17960_/X _18194_/X _24230_/Q _18021_/A VGND VGND VPWR VPWR _24230_/D sky130_fd_sc_hd__o22a_4
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358_ _14355_/X _14357_/Y _12063_/A _14355_/X VGND VGND VPWR VPWR _25148_/D sky130_fd_sc_hd__a2bb2o_4
X_17146_ _16960_/Y _17151_/A VGND VGND VPWR VPWR _17146_/Y sky130_fd_sc_hd__nand2_4
XFILLER_7_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22841__A1 _12228_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24154__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13309_ _13309_/A _13309_/B _13308_/X VGND VGND VPWR VPWR _13309_/X sky130_fd_sc_hd__and3_4
XANTENNA__13468__A _13467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17077_ _17050_/A _17091_/B _17048_/B _17047_/A VGND VGND VPWR VPWR _17077_/X sky130_fd_sc_hd__or4_4
X_14289_ _12027_/D VGND VGND VPWR VPWR _14291_/C sky130_fd_sc_hd__inv_2
X_16028_ _16026_/Y _16022_/X _15959_/X _16027_/X VGND VGND VPWR VPWR _16028_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13334__B2 _11965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14531__B1 _25102_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13187__B _18944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15874__A3 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18273__A1 _13784_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_16_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17979_ _18217_/A _17970_/X _17979_/C VGND VGND VPWR VPWR _17994_/B sky130_fd_sc_hd__or3_4
X_19718_ _19717_/Y _19712_/X _19599_/X _19712_/X VGND VGND VPWR VPWR _23632_/D sky130_fd_sc_hd__a2bb2o_4
X_20990_ _24324_/Q _20990_/B VGND VGND VPWR VPWR _20990_/X sky130_fd_sc_hd__and2_4
XFILLER_81_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16036__B1 _11796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12230__A2_N _12228_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19649_ _19648_/Y _19646_/X _19547_/X _19646_/X VGND VGND VPWR VPWR _19649_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22660_ _22660_/A _22565_/X VGND VGND VPWR VPWR _22662_/B sky130_fd_sc_hd__or2_4
XFILLER_59_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24995__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21611_ _21608_/A _20117_/Y VGND VGND VPWR VPWR _21611_/X sky130_fd_sc_hd__or2_4
XANTENNA__23321__A2 _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20467__C _20481_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22591_ _22476_/X _22590_/X _21285_/A _24818_/Q _22551_/X VGND VGND VPWR VPWR _22591_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17536__B1 _11798_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16019__A _24725_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12245__A2_N _24758_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24924__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24330_ _24330_/CLK _24330_/D HRESETn VGND VGND VPWR VPWR _17199_/A sky130_fd_sc_hd__dfrtp_4
X_21542_ _21542_/A _22111_/B VGND VGND VPWR VPWR _21542_/Y sky130_fd_sc_hd__nand2_4
XFILLER_90_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23140__A _24761_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_16_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15858__A _15852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19289__B1 _19155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24261_ _24689_/CLK _24261_/D HRESETn VGND VGND VPWR VPWR _24261_/Q sky130_fd_sc_hd__dfrtp_4
X_21473_ _21478_/A VGND VGND VPWR VPWR _21670_/A sky130_fd_sc_hd__buf_2
XFILLER_14_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23212_ _23271_/A _23212_/B VGND VGND VPWR VPWR _23222_/B sky130_fd_sc_hd__and2_4
X_20424_ _20423_/X VGND VGND VPWR VPWR _20424_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24192_ _23377_/CLK _24192_/D HRESETn VGND VGND VPWR VPWR _17453_/A sky130_fd_sc_hd__dfrtp_4
X_23143_ _23143_/A _23143_/B VGND VGND VPWR VPWR _23155_/B sky130_fd_sc_hd__and2_4
X_20355_ _21462_/B _20352_/X _19632_/A _20352_/X VGND VGND VPWR VPWR _20355_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15865__A3 _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23074_ _24727_/Q _21021_/X _21050_/X _23073_/X VGND VGND VPWR VPWR _23074_/X sky130_fd_sc_hd__a211o_4
X_20286_ _21915_/B _20283_/X _19985_/X _20283_/X VGND VGND VPWR VPWR _20286_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22596__B1 _25518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22025_ _22025_/A _22023_/X _22025_/C VGND VGND VPWR VPWR _22025_/X sky130_fd_sc_hd__and3_4
XANTENNA__15593__A _15588_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18264__A1 _13795_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19213__B1 _19212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11990_ _11990_/A VGND VGND VPWR VPWR _11990_/Y sky130_fd_sc_hd__inv_2
X_23976_ _23978_/CLK _23976_/D HRESETn VGND VGND VPWR VPWR _20638_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22927_ _22927_/A VGND VGND VPWR VPWR _23171_/B sky130_fd_sc_hd__buf_2
XFILLER_45_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16041__A1_N _16039_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20933__A1_N _20909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13660_ _24039_/Q _13659_/X VGND VGND VPWR VPWR _13661_/B sky130_fd_sc_hd__or2_4
XANTENNA__17313__A _17252_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22858_ _22470_/X _22857_/X _21416_/X _12555_/A _22766_/X VGND VGND VPWR VPWR _22859_/B
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_7_36_0_HCLK clkbuf_6_18_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_73_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12611_ _12670_/A _12611_/B _12666_/A VGND VGND VPWR VPWR _12611_/X sky130_fd_sc_hd__or3_4
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21809_ _21485_/A _21807_/X _21808_/X VGND VGND VPWR VPWR _21809_/X sky130_fd_sc_hd__and3_4
X_13591_ _14620_/B VGND VGND VPWR VPWR _13591_/Y sky130_fd_sc_hd__inv_2
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_99_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_99_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22789_ _23054_/A _22789_/B VGND VGND VPWR VPWR _22789_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24665__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15330_ _24990_/Q _15329_/Y VGND VGND VPWR VPWR _15330_/X sky130_fd_sc_hd__or2_4
XANTENNA__22873__B _22873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12542_ _12542_/A VGND VGND VPWR VPWR _12542_/Y sky130_fd_sc_hd__inv_2
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24528_ _24557_/CLK _16559_/X HRESETn VGND VGND VPWR VPWR _24528_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15261_ _25004_/Q _15261_/B VGND VGND VPWR VPWR _15261_/X sky130_fd_sc_hd__or2_4
XFILLER_32_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15768__A _18254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12473_ _12475_/B VGND VGND VPWR VPWR _12474_/B sky130_fd_sc_hd__inv_2
XANTENNA__23076__A1 _12841_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24459_ _25020_/CLK _24459_/D HRESETn VGND VGND VPWR VPWR _24459_/Q sky130_fd_sc_hd__dfrtp_4
X_14212_ _14212_/A VGND VGND VPWR VPWR _14212_/Y sky130_fd_sc_hd__inv_2
X_17000_ _16017_/Y _17085_/A _16017_/Y _17085_/A VGND VGND VPWR VPWR _17003_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15192_ _15070_/B _15069_/X _15171_/B VGND VGND VPWR VPWR _15193_/B sky130_fd_sc_hd__or3_4
XANTENNA__22823__A1 _12286_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_HCLK clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_3_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12904__B _12903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14143_ _14110_/X _14142_/X _25127_/Q _14136_/X VGND VGND VPWR VPWR _14143_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_10_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14074_ _23994_/Q _14069_/X _14073_/X _14007_/X _14066_/X VGND VGND VPWR VPWR _25226_/D
+ sky130_fd_sc_hd__a32o_4
X_18951_ _18951_/A VGND VGND VPWR VPWR _18951_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13025_ _12999_/X _13017_/D _12306_/Y VGND VGND VPWR VPWR _13025_/X sky130_fd_sc_hd__o21a_4
X_17902_ _17887_/Y _17901_/X _17887_/Y _17901_/X VGND VGND VPWR VPWR _24244_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18882_ _18881_/X VGND VGND VPWR VPWR _18882_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25453__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17833_ _17756_/A _17833_/B VGND VGND VPWR VPWR _17834_/C sky130_fd_sc_hd__or2_4
XANTENNA__19204__B1 _19136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17764_ _17792_/C _17771_/A VGND VGND VPWR VPWR _17765_/D sky130_fd_sc_hd__or2_4
XFILLER_82_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14976_ _14975_/Y _16850_/A _14990_/A _14944_/Y VGND VGND VPWR VPWR _14976_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16018__B1 _11771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19503_ _19502_/Y _19500_/X _11943_/X _19500_/X VGND VGND VPWR VPWR _19503_/X sky130_fd_sc_hd__a2bb2o_4
X_16715_ _21582_/A _16712_/X _16442_/X _16712_/X VGND VGND VPWR VPWR _24468_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13927_ _13927_/A _13927_/B _13895_/A _13927_/D VGND VGND VPWR VPWR _13946_/D sky130_fd_sc_hd__or4_4
X_17695_ _17695_/A VGND VGND VPWR VPWR _17696_/B sky130_fd_sc_hd__inv_2
XFILLER_19_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18319__A _17700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19434_ _19433_/Y _19431_/X _19364_/X _19431_/X VGND VGND VPWR VPWR _23729_/D sky130_fd_sc_hd__a2bb2o_4
X_16646_ _16658_/A VGND VGND VPWR VPWR _16646_/X sky130_fd_sc_hd__buf_2
XFILLER_35_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13858_ _13851_/X VGND VGND VPWR VPWR _13858_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12809_ _12887_/A _24795_/Q _12887_/A _24795_/Q VGND VGND VPWR VPWR _12815_/B sky130_fd_sc_hd__a2bb2o_4
X_19365_ _19363_/Y _19361_/X _19364_/X _19361_/X VGND VGND VPWR VPWR _23753_/D sky130_fd_sc_hd__a2bb2o_4
X_16577_ _24520_/Q VGND VGND VPWR VPWR _16577_/Y sky130_fd_sc_hd__inv_2
X_13789_ _15662_/A _13789_/B _12095_/Y _13789_/D VGND VGND VPWR VPWR _21027_/B sky130_fd_sc_hd__or4_4
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18316_ _18298_/X _18301_/B _18295_/Y VGND VGND VPWR VPWR _18316_/X sky130_fd_sc_hd__o21a_4
XFILLER_15_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15528_ _24919_/Q VGND VGND VPWR VPWR _15528_/Y sky130_fd_sc_hd__inv_2
X_19296_ _19293_/Y _19288_/X _19294_/X _19295_/X VGND VGND VPWR VPWR _19296_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21865__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24335__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18247_ HWDATA[7] VGND VGND VPWR VPWR _18247_/X sky130_fd_sc_hd__buf_2
X_15459_ _13893_/B _20602_/A _15446_/A _13927_/A _15434_/X VGND VGND VPWR VPWR _15459_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_129_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14902__A2_N _14900_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18178_ _17928_/A _18178_/B _18178_/C VGND VGND VPWR VPWR _18178_/X sky130_fd_sc_hd__and3_4
XFILLER_89_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17129_ _17044_/B _17128_/X VGND VGND VPWR VPWR _17130_/B sky130_fd_sc_hd__or2_4
XFILLER_85_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20140_ _20140_/A VGND VGND VPWR VPWR _20140_/X sky130_fd_sc_hd__buf_2
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22578__B1 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23970__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20071_ _20064_/X _18325_/X _18254_/X _13348_/B _20066_/X VGND VGND VPWR VPWR _23504_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_131_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19443__B1 _19420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25194__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12830__A _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16257__B1 _16064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22593__A3 _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23830_ _25054_/CLK _19147_/X VGND VGND VPWR VPWR _23830_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16272__A3 _16270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21862__B _21862_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23761_ _23828_/CLK _23761_/D VGND VGND VPWR VPWR _18083_/B sky130_fd_sc_hd__dfxtp_4
X_20973_ _24108_/Q _24106_/Q _24107_/Q _20972_/X VGND VGND VPWR VPWR _20973_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17133__A _17038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25500_ _25497_/CLK _11915_/X HRESETn VGND VGND VPWR VPWR _11877_/A sky130_fd_sc_hd__dfrtp_4
X_22712_ _22266_/X VGND VGND VPWR VPWR _22712_/X sky130_fd_sc_hd__buf_2
X_23692_ _23384_/CLK _19540_/X VGND VGND VPWR VPWR _22386_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_41_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25431_ _25449_/CLK _12476_/X HRESETn VGND VGND VPWR VPWR _12474_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22643_ _22611_/X _22618_/Y _22622_/X _22642_/Y VGND VGND VPWR VPWR HRDATA[12] sky130_fd_sc_hd__or4_4
XANTENNA__17509__B1 _11828_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12277__A _12277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25362_ _25330_/CLK _12962_/X HRESETn VGND VGND VPWR VPWR _25362_/Q sky130_fd_sc_hd__dfrtp_4
X_22574_ _22574_/A _22571_/X _22574_/C VGND VGND VPWR VPWR _22574_/X sky130_fd_sc_hd__and3_4
XFILLER_55_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24313_ _24883_/CLK _24313_/D HRESETn VGND VGND VPWR VPWR _17436_/A sky130_fd_sc_hd__dfrtp_4
X_21525_ _21525_/A VGND VGND VPWR VPWR _22879_/A sky130_fd_sc_hd__buf_2
XFILLER_107_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15588__A _15588_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25293_ _25478_/CLK _25293_/D HRESETn VGND VGND VPWR VPWR _25293_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14492__A _25101_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24005__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24244_ _24186_/CLK _24244_/D HRESETn VGND VGND VPWR VPWR _24244_/Q sky130_fd_sc_hd__dfrtp_4
X_21456_ _21456_/A _19882_/Y VGND VGND VPWR VPWR _21460_/B sky130_fd_sc_hd__or2_4
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20407_ _23375_/Q VGND VGND VPWR VPWR _20407_/Y sky130_fd_sc_hd__inv_2
X_24175_ _24171_/CLK _18489_/Y HRESETn VGND VGND VPWR VPWR _18455_/A sky130_fd_sc_hd__dfrtp_4
X_21387_ _21383_/X _21386_/X _14676_/A VGND VGND VPWR VPWR _21387_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16496__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23126_ _23126_/A VGND VGND VPWR VPWR _23128_/A sky130_fd_sc_hd__buf_2
X_20338_ _20338_/A _20338_/B _19888_/C VGND VGND VPWR VPWR _20338_/X sky130_fd_sc_hd__or3_4
XANTENNA__15838__A3 _15768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19434__B1 _19364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17308__A _17252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23057_ _22520_/A VGND VGND VPWR VPWR _23057_/X sky130_fd_sc_hd__buf_2
X_20269_ _20268_/Y _20266_/X _19797_/A _20266_/X VGND VGND VPWR VPWR _23430_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16248__B1 _16143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22008_ _22016_/A _19872_/Y VGND VGND VPWR VPWR _22011_/B sky130_fd_sc_hd__or2_4
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14830_ _14825_/X _14829_/X _25042_/Q _14825_/X VGND VGND VPWR VPWR _14830_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11973_ _21504_/A _11972_/X _11958_/X _13678_/B VGND VGND VPWR VPWR _11976_/A sky130_fd_sc_hd__o22a_4
X_14761_ _14770_/B VGND VGND VPWR VPWR _14772_/A sky130_fd_sc_hd__inv_2
XFILLER_99_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23959_ _23959_/CLK _23959_/D HRESETn VGND VGND VPWR VPWR _20530_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__18139__A _18024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21544__B2 _17416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22741__B1 _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24846__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16500_ _16497_/Y _16499_/X _16325_/X _16499_/X VGND VGND VPWR VPWR _16500_/X sky130_fd_sc_hd__a2bb2o_4
X_13712_ _13689_/A _13689_/B VGND VGND VPWR VPWR _13712_/Y sky130_fd_sc_hd__nand2_4
X_14692_ _21391_/A VGND VGND VPWR VPWR _14693_/A sky130_fd_sc_hd__buf_2
X_17480_ _24310_/Q VGND VGND VPWR VPWR _17480_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16420__B1 _16231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16431_ _15099_/Y _16429_/X _16147_/X _16429_/X VGND VGND VPWR VPWR _16431_/X sky130_fd_sc_hd__a2bb2o_4
X_13643_ _13536_/Y _13643_/B VGND VGND VPWR VPWR _13644_/A sky130_fd_sc_hd__or2_4
XFILLER_38_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20887__A1_N _20882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19150_ _19148_/Y _19144_/X _19149_/X _19130_/A VGND VGND VPWR VPWR _19150_/X sky130_fd_sc_hd__a2bb2o_4
X_13574_ _25245_/Q _13573_/A _13572_/Y _13573_/Y VGND VGND VPWR VPWR _13574_/X sky130_fd_sc_hd__o22a_4
X_16362_ _16361_/Y _16356_/X _15986_/X _16356_/X VGND VGND VPWR VPWR _24601_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21847__A2 _13496_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18101_ _18133_/A _18101_/B VGND VGND VPWR VPWR _18101_/X sky130_fd_sc_hd__or2_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _25398_/Q _12523_/Y _12524_/Y _24868_/Q VGND VGND VPWR VPWR _12525_/X sky130_fd_sc_hd__a2bb2o_4
X_15313_ _15313_/A _15313_/B VGND VGND VPWR VPWR _15314_/C sky130_fd_sc_hd__or2_4
X_16293_ _24626_/Q VGND VGND VPWR VPWR _16293_/Y sky130_fd_sc_hd__inv_2
X_19081_ _23853_/Q VGND VGND VPWR VPWR _19081_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_123_0_HCLK clkbuf_7_61_0_HCLK/X VGND VGND VPWR VPWR _24581_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18032_ _18217_/A _18027_/X _18032_/C VGND VGND VPWR VPWR _18040_/B sky130_fd_sc_hd__or3_4
Xclkbuf_8_186_0_HCLK clkbuf_7_93_0_HCLK/X VGND VGND VPWR VPWR _23398_/CLK sky130_fd_sc_hd__clkbuf_1
X_12456_ _12429_/X _12454_/X _12456_/C VGND VGND VPWR VPWR _25435_/D sky130_fd_sc_hd__and3_4
X_15244_ _15239_/A _15239_/B _15199_/X _15240_/Y VGND VGND VPWR VPWR _15245_/A sky130_fd_sc_hd__a211o_4
XANTENNA__20810__A1_N _20680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15175_ _15166_/C _15173_/X _15174_/X _15167_/Y VGND VGND VPWR VPWR _15176_/A sky130_fd_sc_hd__a211o_4
X_12387_ _25451_/Q _12387_/B VGND VGND VPWR VPWR _12389_/B sky130_fd_sc_hd__or2_4
XFILLER_67_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14126_ _14108_/X VGND VGND VPWR VPWR _14132_/A sky130_fd_sc_hd__buf_2
XANTENNA__16487__B1 _16401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19983_ _22029_/B _19974_/X _19981_/X _19982_/X VGND VGND VPWR VPWR _19983_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14057_ _14078_/A VGND VGND VPWR VPWR _14057_/X sky130_fd_sc_hd__buf_2
X_18934_ _13347_/B VGND VGND VPWR VPWR _18934_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12650__A _12665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16239__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13008_ _13002_/B _13008_/B VGND VGND VPWR VPWR _13017_/D sky130_fd_sc_hd__and2_4
XFILLER_132_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18865_ _18849_/X _18865_/B _18865_/C _18865_/D VGND VGND VPWR VPWR _18865_/X sky130_fd_sc_hd__or4_4
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17816_ _16941_/Y _17810_/X _17780_/X _17813_/B VGND VGND VPWR VPWR _17817_/A sky130_fd_sc_hd__a211o_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18796_ _18796_/A VGND VGND VPWR VPWR _18796_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17747_ _17744_/Y _16928_/Y _17747_/C _17747_/D VGND VGND VPWR VPWR _17747_/X sky130_fd_sc_hd__or4_4
XFILLER_36_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14959_ _15219_/B _24418_/Q _14903_/X _14904_/Y VGND VGND VPWR VPWR _14963_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13473__B1 _13472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18049__A _18177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24587__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17678_ _17512_/Y _17665_/X VGND VGND VPWR VPWR _17679_/C sky130_fd_sc_hd__nand2_4
XANTENNA__22794__A _22794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24516__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16411__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19417_ _18171_/B VGND VGND VPWR VPWR _19417_/Y sky130_fd_sc_hd__inv_2
X_16629_ _13741_/A VGND VGND VPWR VPWR _16629_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17888__A _17700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12097__A _12096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_2_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19348_ _19348_/A VGND VGND VPWR VPWR _19348_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21838__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_82_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_82_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19279_ _21607_/B _19278_/X _16885_/X _19278_/X VGND VGND VPWR VPWR _23783_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12825__A _25375_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21310_ _15671_/A VGND VGND VPWR VPWR _22927_/A sky130_fd_sc_hd__buf_2
XFILLER_11_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22290_ _22289_/Y _22278_/X _13128_/A _21278_/X VGND VGND VPWR VPWR _22290_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22799__B1 _22798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21241_ _21240_/X _20122_/Y VGND VGND VPWR VPWR _21241_/X sky130_fd_sc_hd__or2_4
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21857__B _23082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25375__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20274__A1 _23428_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21172_ _21184_/A _19487_/Y VGND VGND VPWR VPWR _21172_/X sky130_fd_sc_hd__or2_4
XANTENNA__25304__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20123_ _19841_/A VGND VGND VPWR VPWR _20123_/X sky130_fd_sc_hd__buf_2
XANTENNA__19416__B1 _19370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20054_ _23512_/Q VGND VGND VPWR VPWR _20054_/Y sky130_fd_sc_hd__inv_2
X_24931_ _23711_/CLK _15500_/X HRESETn VGND VGND VPWR VPWR _11727_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_112_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24862_ _24457_/CLK _15734_/X HRESETn VGND VGND VPWR VPWR _24862_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_61_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23813_ _23832_/CLK _19194_/X VGND VGND VPWR VPWR _19193_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12267__B2 _24765_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13464__B1 _25313_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24793_ _24800_/CLK _15880_/X HRESETn VGND VGND VPWR VPWR _22967_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14487__A _25103_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ _23446_/CLK _19390_/X VGND VGND VPWR VPWR _18101_/B sky130_fd_sc_hd__dfxtp_4
X_20956_ _12010_/A _20958_/B VGND VGND VPWR VPWR _20956_/X sky130_fd_sc_hd__and2_4
XANTENNA__15205__A1 _15069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24257__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16402__B1 _16401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_5_31_0_HCLK_A clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _23384_/CLK _19591_/X VGND VGND VPWR VPWR _22220_/A sky130_fd_sc_hd__dfxtp_4
X_20887_ _20882_/X _20885_/Y _16682_/A _20886_/X VGND VGND VPWR VPWR _24044_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25414_ _25411_/CLK _25414_/D HRESETn VGND VGND VPWR VPWR _12524_/A sky130_fd_sc_hd__dfrtp_4
X_22626_ _24747_/Q _22626_/B VGND VGND VPWR VPWR _22626_/X sky130_fd_sc_hd__or2_4
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25345_ _23370_/CLK _25345_/D HRESETn VGND VGND VPWR VPWR _25345_/Q sky130_fd_sc_hd__dfrtp_4
X_22557_ _21582_/B VGND VGND VPWR VPWR _22922_/A sky130_fd_sc_hd__buf_2
X_12310_ _25343_/Q _12308_/Y _25349_/Q _12309_/Y VGND VGND VPWR VPWR _12313_/C sky130_fd_sc_hd__a2bb2o_4
X_21508_ _21507_/Y VGND VGND VPWR VPWR _22035_/A sky130_fd_sc_hd__buf_2
X_13290_ _13251_/A _19757_/A VGND VGND VPWR VPWR _13290_/X sky130_fd_sc_hd__or2_4
X_25276_ _25279_/CLK _25276_/D HRESETn VGND VGND VPWR VPWR _11685_/A sky130_fd_sc_hd__dfrtp_4
X_22488_ _22778_/A _22488_/B _22488_/C _22487_/X VGND VGND VPWR VPWR _22488_/X sky130_fd_sc_hd__or4_4
X_12241_ _12462_/A VGND VGND VPWR VPWR _12242_/A sky130_fd_sc_hd__inv_2
X_24227_ _24715_/CLK _24227_/D HRESETn VGND VGND VPWR VPWR _24227_/Q sky130_fd_sc_hd__dfrtp_4
X_21439_ _11720_/B VGND VGND VPWR VPWR _22821_/A sky130_fd_sc_hd__buf_2
XFILLER_108_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12172_ _13533_/A _12060_/B _15652_/D _13533_/D VGND VGND VPWR VPWR _12173_/A sky130_fd_sc_hd__or4_4
X_24158_ _24159_/CLK _18555_/X HRESETn VGND VGND VPWR VPWR _18467_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25045__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23109_ _23108_/X VGND VGND VPWR VPWR _23109_/Y sky130_fd_sc_hd__inv_2
X_16980_ _16973_/X _16980_/B _16977_/X _16980_/D VGND VGND VPWR VPWR _16990_/C sky130_fd_sc_hd__or4_4
X_24089_ _24089_/CLK _24089_/D HRESETn VGND VGND VPWR VPWR _11994_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_77_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22879__A _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15931_ _15931_/A _15931_/B VGND VGND VPWR VPWR _15967_/A sky130_fd_sc_hd__or2_4
XFILLER_77_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18650_ _24128_/Q VGND VGND VPWR VPWR _18767_/A sky130_fd_sc_hd__buf_2
X_15862_ _15702_/A _15931_/B VGND VGND VPWR VPWR _15863_/A sky130_fd_sc_hd__or2_4
X_17601_ _17885_/B VGND VGND VPWR VPWR _17601_/X sky130_fd_sc_hd__buf_2
X_14813_ _14870_/B _14798_/X _14813_/C VGND VGND VPWR VPWR _14813_/X sky130_fd_sc_hd__or3_4
X_18581_ _18581_/A _18581_/B VGND VGND VPWR VPWR _18582_/B sky130_fd_sc_hd__or2_4
X_15793_ _15793_/A VGND VGND VPWR VPWR _15793_/X sky130_fd_sc_hd__buf_2
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24680__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17532_ _17526_/X _17529_/X _17530_/X _17531_/X VGND VGND VPWR VPWR _17532_/X sky130_fd_sc_hd__or4_4
X_14744_ _21781_/A _14703_/A _14705_/B VGND VGND VPWR VPWR _14744_/X sky130_fd_sc_hd__o21a_4
X_11956_ _11954_/Y _11947_/X _11955_/X _11947_/A VGND VGND VPWR VPWR _11956_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12629__B _12602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17463_ _17462_/Y VGND VGND VPWR VPWR _17472_/A sky130_fd_sc_hd__buf_2
XFILLER_60_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11887_ _11924_/A _11899_/A _11872_/X _11882_/X _11886_/Y VGND VGND VPWR VPWR _11887_/X
+ sky130_fd_sc_hd__a2111o_4
X_14675_ _24936_/Q _11709_/B _14675_/C _13593_/X VGND VGND VPWR VPWR _14675_/X sky130_fd_sc_hd__or4_4
X_19202_ _18056_/B VGND VGND VPWR VPWR _19202_/Y sky130_fd_sc_hd__inv_2
X_16414_ _16433_/A VGND VGND VPWR VPWR _16414_/X sky130_fd_sc_hd__buf_2
X_13626_ _19152_/D _13626_/B VGND VGND VPWR VPWR _13626_/X sky130_fd_sc_hd__and2_4
X_17394_ _20638_/A _20638_/B VGND VGND VPWR VPWR _20642_/B sky130_fd_sc_hd__or2_4
XFILLER_9_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11769__B1 _11767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19133_ _19642_/A VGND VGND VPWR VPWR _19133_/X sky130_fd_sc_hd__buf_2
X_16345_ _16345_/A VGND VGND VPWR VPWR _16345_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13557_ _13557_/A VGND VGND VPWR VPWR _13557_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12508_ _21065_/A _13026_/A VGND VGND VPWR VPWR _12509_/C sky130_fd_sc_hd__or2_4
X_19064_ _19060_/Y _19063_/X _19018_/X _19063_/X VGND VGND VPWR VPWR _19064_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12981__A2 _12866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13488_ _13488_/A VGND VGND VPWR VPWR _13488_/Y sky130_fd_sc_hd__inv_2
X_16276_ _22671_/A _16276_/B VGND VGND VPWR VPWR _16276_/X sky130_fd_sc_hd__or2_4
X_18015_ _18056_/A _19200_/A VGND VGND VPWR VPWR _18015_/X sky130_fd_sc_hd__or2_4
X_12439_ _12438_/X VGND VGND VPWR VPWR _25440_/D sky130_fd_sc_hd__inv_2
X_15227_ _15227_/A _15227_/B VGND VGND VPWR VPWR _15228_/C sky130_fd_sc_hd__or2_4
XFILLER_86_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15158_ _24969_/Q VGND VGND VPWR VPWR _15406_/A sky130_fd_sc_hd__inv_2
XANTENNA__15675__B _15674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14109_ _14108_/X VGND VGND VPWR VPWR _14129_/A sky130_fd_sc_hd__inv_2
XFILLER_102_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13476__A _13475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15089_ _15089_/A VGND VGND VPWR VPWR _15089_/Y sky130_fd_sc_hd__inv_2
X_19966_ _23542_/Q VGND VGND VPWR VPWR _19966_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18917_ _21384_/B _18914_/X _16888_/X _18914_/X VGND VGND VPWR VPWR _18917_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22548__A3 _22127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21693__A _23314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19897_ _19897_/A VGND VGND VPWR VPWR _21937_/B sky130_fd_sc_hd__inv_2
XFILLER_68_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16787__A _16786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24768__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18848_ _24551_/Q _18757_/A _16513_/Y _24123_/Q VGND VGND VPWR VPWR _18849_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18779_ _18778_/X VGND VGND VPWR VPWR _24125_/D sky130_fd_sc_hd__inv_2
X_20810_ _20680_/X _20809_/X _15559_/A _20725_/X VGND VGND VPWR VPWR _20810_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21790_ _21485_/A _21788_/X _21789_/X VGND VGND VPWR VPWR _21790_/X sky130_fd_sc_hd__and3_4
XANTENNA__24350__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20741_ _20738_/Y _20739_/Y _20740_/X VGND VGND VPWR VPWR _20741_/X sky130_fd_sc_hd__o21a_4
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19825__A2_N _19824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23460_ _23434_/CLK _23460_/D VGND VGND VPWR VPWR _23460_/Q sky130_fd_sc_hd__dfxtp_4
X_20672_ _20487_/A _20479_/C _20602_/X VGND VGND VPWR VPWR _20672_/X sky130_fd_sc_hd__o21a_4
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22411_ _21413_/X _22410_/X _22396_/C _12542_/A _22540_/A VGND VGND VPWR VPWR _22411_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12421__A1 _12277_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23391_ _23682_/CLK _23391_/D VGND VGND VPWR VPWR _23391_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12555__A _12555_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15539__A2_N _15535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25130_ _25093_/CLK _25130_/D HRESETn VGND VGND VPWR VPWR _14416_/A sky130_fd_sc_hd__dfstp_4
X_22342_ _21929_/A _22342_/B VGND VGND VPWR VPWR _22342_/X sky130_fd_sc_hd__or2_4
X_25061_ _25044_/CLK _14666_/Y HRESETn VGND VGND VPWR VPWR _25061_/Q sky130_fd_sc_hd__dfrtp_4
X_22273_ _22273_/A _22272_/X VGND VGND VPWR VPWR _22273_/X sky130_fd_sc_hd__or2_4
XANTENNA__12185__B1 _12277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_26_0_HCLK clkbuf_8_27_0_HCLK/A VGND VGND VPWR VPWR _25301_/CLK sky130_fd_sc_hd__clkbuf_1
X_24012_ _24909_/CLK _24012_/D HRESETn VGND VGND VPWR VPWR _24012_/Q sky130_fd_sc_hd__dfrtp_4
X_21224_ _21372_/A VGND VGND VPWR VPWR _21249_/A sky130_fd_sc_hd__buf_2
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_89_0_HCLK clkbuf_8_89_0_HCLK/A VGND VGND VPWR VPWR _23989_/CLK sky130_fd_sc_hd__clkbuf_1
X_21155_ _15336_/A _15852_/A _21314_/B VGND VGND VPWR VPWR _21155_/X sky130_fd_sc_hd__and3_4
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12290__A _12290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20106_ _20105_/X VGND VGND VPWR VPWR _20106_/X sky130_fd_sc_hd__buf_2
X_21086_ _24599_/Q _22587_/B VGND VGND VPWR VPWR _21086_/X sky130_fd_sc_hd__or2_4
X_20037_ _20035_/Y _20036_/X _19992_/X _20036_/X VGND VGND VPWR VPWR _20037_/X sky130_fd_sc_hd__a2bb2o_4
X_24914_ _25255_/CLK _24914_/D HRESETn VGND VGND VPWR VPWR _24914_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23307__B _21519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24438__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16623__B1 _16366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21108__A _15638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24845_ _24842_/CLK _15769_/X HRESETn VGND VGND VPWR VPWR _24845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11810_ _11807_/Y _11805_/X _11809_/X _11805_/X VGND VGND VPWR VPWR _11810_/X sky130_fd_sc_hd__a2bb2o_4
X_12790_ _12780_/X _12783_/X _12790_/C _12789_/X VGND VGND VPWR VPWR _12790_/X sky130_fd_sc_hd__or4_4
X_21988_ _24243_/Q _20331_/Y _21985_/X _21987_/X VGND VGND VPWR VPWR _21989_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24091__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24776_ _24821_/CLK _15906_/X HRESETn VGND VGND VPWR VPWR _24776_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17179__B2 _17178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11750_/A VGND VGND VPWR VPWR _11741_/X sky130_fd_sc_hd__buf_2
XFILLER_26_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20939_ _20939_/A _20939_/B VGND VGND VPWR VPWR _20939_/X sky130_fd_sc_hd__and2_4
XFILLER_15_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20183__B1 _20096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23727_ _23722_/CLK _19439_/X VGND VGND VPWR VPWR _18140_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24020__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _13676_/A _11664_/Y _25279_/Q _11671_/Y VGND VGND VPWR VPWR _11675_/C sky130_fd_sc_hd__a2bb2o_4
X_14460_ _14458_/Y _14454_/X _14418_/X _14459_/X VGND VGND VPWR VPWR _25114_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23658_ _24197_/CLK _23658_/D VGND VGND VPWR VPWR _23658_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13411_ _13379_/A _13411_/B VGND VGND VPWR VPWR _13411_/X sky130_fd_sc_hd__or2_4
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ _16355_/A VGND VGND VPWR VPWR _14391_/X sky130_fd_sc_hd__buf_2
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22609_ _24445_/Q _22525_/X _22526_/X VGND VGND VPWR VPWR _22609_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25297__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23589_ _24089_/CLK _23589_/D VGND VGND VPWR VPWR _23589_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13342_ _13301_/X _13340_/X _13341_/X VGND VGND VPWR VPWR _13342_/X sky130_fd_sc_hd__and3_4
X_16130_ _16130_/A VGND VGND VPWR VPWR _16130_/Y sky130_fd_sc_hd__inv_2
X_25328_ _24836_/CLK _25328_/D HRESETn VGND VGND VPWR VPWR _12377_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15049__A1_N _14888_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25226__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13273_ _13417_/A _13273_/B VGND VGND VPWR VPWR _13274_/C sky130_fd_sc_hd__or2_4
X_16061_ _15623_/A VGND VGND VPWR VPWR _16061_/X sky130_fd_sc_hd__buf_2
X_25259_ _25070_/CLK _25259_/D HRESETn VGND VGND VPWR VPWR _25259_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18152__A _18184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12176__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12224_ _21526_/A VGND VGND VPWR VPWR _12224_/Y sky130_fd_sc_hd__inv_2
X_15012_ _15004_/X _15012_/B _15012_/C _15012_/D VGND VGND VPWR VPWR _15012_/X sky130_fd_sc_hd__or4_4
XANTENNA__21435__B1 _24808_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19820_ _19819_/Y _19815_/X _19771_/X _19802_/Y VGND VGND VPWR VPWR _19820_/X sky130_fd_sc_hd__a2bb2o_4
X_12155_ _12151_/A _12148_/A _12153_/Y VGND VGND VPWR VPWR _12155_/X sky130_fd_sc_hd__o21a_4
XFILLER_97_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11809__A _11809_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23188__B1 _11756_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19751_ _19750_/X VGND VGND VPWR VPWR _19751_/Y sky130_fd_sc_hd__inv_2
X_12086_ _12073_/Y VGND VGND VPWR VPWR _12086_/X sky130_fd_sc_hd__buf_2
X_16963_ _16958_/X _16959_/X _16961_/X _16962_/X VGND VGND VPWR VPWR _16990_/A sky130_fd_sc_hd__or4_4
XANTENNA__24861__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18702_ _18738_/A _18700_/X _18701_/Y VGND VGND VPWR VPWR _24144_/D sky130_fd_sc_hd__and3_4
X_15914_ _15912_/X VGND VGND VPWR VPWR _15915_/B sky130_fd_sc_hd__inv_2
X_19682_ _23644_/Q VGND VGND VPWR VPWR _19682_/Y sky130_fd_sc_hd__inv_2
X_16894_ _16103_/Y _17742_/A _16103_/Y _17742_/A VGND VGND VPWR VPWR _16895_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22121__B _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18633_ _18633_/A VGND VGND VPWR VPWR _18682_/B sky130_fd_sc_hd__inv_2
X_15845_ _15845_/A VGND VGND VPWR VPWR _15845_/X sky130_fd_sc_hd__buf_2
XFILLER_94_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18564_ _18469_/B _18576_/B VGND VGND VPWR VPWR _18574_/B sky130_fd_sc_hd__or2_4
X_15776_ _15552_/Y _15646_/X _15774_/X _24841_/Q _15775_/X VGND VGND VPWR VPWR _15776_/X
+ sky130_fd_sc_hd__a32o_4
X_12988_ _12988_/A _13057_/A _12358_/Y _12349_/Y VGND VGND VPWR VPWR _12989_/C sky130_fd_sc_hd__or4_4
XFILLER_73_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17515_ _17515_/A VGND VGND VPWR VPWR _17597_/A sky130_fd_sc_hd__inv_2
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14727_ _22036_/A VGND VGND VPWR VPWR _14727_/Y sky130_fd_sc_hd__inv_2
X_11939_ _19618_/A VGND VGND VPWR VPWR _11939_/X sky130_fd_sc_hd__buf_2
X_18495_ _18517_/A _18495_/B _18494_/X VGND VGND VPWR VPWR _24174_/D sky130_fd_sc_hd__and3_4
XANTENNA__16917__B2 _16916_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17170__A1_N _22273_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12583__A2_N _24846_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17446_ _14675_/C VGND VGND VPWR VPWR _17700_/C sky130_fd_sc_hd__buf_2
X_14658_ _14658_/A _13619_/X VGND VGND VPWR VPWR _14659_/B sky130_fd_sc_hd__or2_4
X_13609_ _18987_/D _13609_/B VGND VGND VPWR VPWR _13609_/X sky130_fd_sc_hd__and2_4
XANTENNA__12403__A1 _12385_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17377_ _17199_/Y _17377_/B VGND VGND VPWR VPWR _17381_/B sky130_fd_sc_hd__or2_4
X_14589_ _14570_/A _14570_/B VGND VGND VPWR VPWR _14589_/X sky130_fd_sc_hd__or2_4
XANTENNA__25131__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19116_ _13338_/B VGND VGND VPWR VPWR _19116_/Y sky130_fd_sc_hd__inv_2
X_16328_ _16327_/Y _16324_/X _16228_/X _16324_/X VGND VGND VPWR VPWR _16328_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17885__B _17885_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17342__A1 _17249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16899__A2_N _16898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19047_ _19047_/A VGND VGND VPWR VPWR _19047_/Y sky130_fd_sc_hd__inv_2
X_16259_ _16192_/A VGND VGND VPWR VPWR _16259_/X sky130_fd_sc_hd__buf_2
XANTENNA__18062__A _13610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_242_0_HCLK clkbuf_8_243_0_HCLK/A VGND VGND VPWR VPWR _24868_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18997__A _18996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24949__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16853__B1 _16852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19949_ _19949_/A VGND VGND VPWR VPWR _19949_/Y sky130_fd_sc_hd__inv_2
X_22960_ _22955_/Y _22959_/Y _22850_/X VGND VGND VPWR VPWR _22961_/D sky130_fd_sc_hd__o21a_4
XANTENNA__24531__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16605__B1 _16604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21911_ _21895_/X _21910_/X _21270_/X VGND VGND VPWR VPWR _21911_/X sky130_fd_sc_hd__a21o_4
XFILLER_55_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22891_ _22464_/A VGND VGND VPWR VPWR _23140_/B sky130_fd_sc_hd__buf_2
XANTENNA__20952__A2 _14620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21842_ _14421_/Y _14223_/A _14444_/Y _22316_/B VGND VGND VPWR VPWR _21842_/X sky130_fd_sc_hd__o22a_4
XFILLER_23_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24630_ _24612_/CLK _24630_/D HRESETn VGND VGND VPWR VPWR _24630_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24561_ _24561_/CLK _16472_/X HRESETn VGND VGND VPWR VPWR _24561_/Q sky130_fd_sc_hd__dfrtp_4
X_21773_ _21630_/A _20091_/Y VGND VGND VPWR VPWR _21774_/C sky130_fd_sc_hd__or2_4
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20724_ _20724_/A VGND VGND VPWR VPWR _20747_/A sky130_fd_sc_hd__inv_2
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23512_ _25264_/CLK _23512_/D VGND VGND VPWR VPWR _23512_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24492_ _24492_/CLK _16656_/X HRESETn VGND VGND VPWR VPWR _24492_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23103__B1 _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23443_ _25316_/CLK _23443_/D VGND VGND VPWR VPWR _13214_/B sky130_fd_sc_hd__dfxtp_4
X_20655_ _17399_/B VGND VGND VPWR VPWR _20655_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22457__A2 _23126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25390__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_52_0_HCLK clkbuf_6_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23374_ _24187_/CLK _23374_/D VGND VGND VPWR VPWR _23374_/Q sky130_fd_sc_hd__dfxtp_4
X_20586_ _23943_/Q _18880_/X _18882_/Y VGND VGND VPWR VPWR _20586_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_87_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22325_ _17717_/A _22325_/B VGND VGND VPWR VPWR _22325_/X sky130_fd_sc_hd__or2_4
X_25113_ _25113_/CLK _14462_/X HRESETn VGND VGND VPWR VPWR _25113_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19068__A _19062_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15895__B2 _15864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25044_ _25044_/CLK _25044_/D HRESETn VGND VGND VPWR VPWR _13598_/C sky130_fd_sc_hd__dfrtp_4
X_22256_ _21681_/A _22248_/X _22255_/X VGND VGND VPWR VPWR _22256_/X sky130_fd_sc_hd__and3_4
XFILLER_133_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20007__A _20014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21207_ _21160_/X _21197_/X _21207_/C VGND VGND VPWR VPWR _21207_/X sky130_fd_sc_hd__or3_4
X_22187_ _22153_/X _22157_/X _22179_/X _22187_/D VGND VGND VPWR VPWR _22293_/A sky130_fd_sc_hd__or4_4
XFILLER_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24619__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21138_ _13789_/D _21130_/X _12066_/X _21137_/X VGND VGND VPWR VPWR _21138_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13960_ _13960_/A VGND VGND VPWR VPWR _13960_/Y sky130_fd_sc_hd__inv_2
X_21069_ _21069_/A VGND VGND VPWR VPWR _23019_/B sky130_fd_sc_hd__buf_2
XFILLER_47_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24272__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12911_ _12911_/A VGND VGND VPWR VPWR _12911_/Y sky130_fd_sc_hd__inv_2
X_13891_ _13926_/C _24958_/Q _13958_/D VGND VGND VPWR VPWR _13892_/A sky130_fd_sc_hd__or3_4
XFILLER_19_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24201__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15630_ _15629_/Y _15626_/X _15471_/X _15626_/X VGND VGND VPWR VPWR _24884_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12842_ _12842_/A _12959_/A _12819_/A _12761_/Y VGND VGND VPWR VPWR _12842_/X sky130_fd_sc_hd__or4_4
X_24828_ _24868_/CLK _24828_/D HRESETn VGND VGND VPWR VPWR _12308_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22145__A1 _15708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20677__A _20676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22145__B2 _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15561_ _15580_/A VGND VGND VPWR VPWR _15561_/X sky130_fd_sc_hd__buf_2
XFILLER_76_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12773_ _12771_/A _12772_/A _12841_/B _12772_/Y VGND VGND VPWR VPWR _12773_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22696__A2 _22406_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25478__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24759_ _24759_/CLK _24759_/D HRESETn VGND VGND VPWR VPWR _12207_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13830__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14675__A _24936_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17291_/X VGND VGND VPWR VPWR _17304_/B sky130_fd_sc_hd__inv_2
XPHY_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _20441_/B VGND VGND VPWR VPWR _14512_/Y sky130_fd_sc_hd__inv_2
X_11724_ _12068_/A _11723_/Y VGND VGND VPWR VPWR _11725_/B sky130_fd_sc_hd__or2_4
X_18280_ _18280_/A VGND VGND VPWR VPWR _18280_/X sky130_fd_sc_hd__buf_2
XPHY_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _11707_/Y _15491_/X HWRITE _15491_/X VGND VGND VPWR VPWR _24936_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25407__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22892__A _22892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17202_/X _17231_/B VGND VGND VPWR VPWR _17231_/X sky130_fd_sc_hd__or2_4
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11655_/A VGND VGND VPWR VPWR _11701_/B sky130_fd_sc_hd__inv_2
X_14443_ _14441_/Y _14437_/X _14418_/X _14442_/X VGND VGND VPWR VPWR _25122_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17162_ _17162_/A _17162_/B VGND VGND VPWR VPWR _17163_/B sky130_fd_sc_hd__or2_4
XFILLER_7_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22177__A1_N _20500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14374_ _14373_/Y VGND VGND VPWR VPWR _20496_/C sky130_fd_sc_hd__buf_2
XANTENNA__25060__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16113_ _16094_/A VGND VGND VPWR VPWR _16113_/X sky130_fd_sc_hd__buf_2
XANTENNA__21301__A _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13325_ _13392_/A _13325_/B VGND VGND VPWR VPWR _13325_/X sky130_fd_sc_hd__or2_4
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17093_ _17007_/Y _17092_/X VGND VGND VPWR VPWR _17093_/X sky130_fd_sc_hd__or2_4
X_16044_ _16044_/A VGND VGND VPWR VPWR _16044_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13256_ _13366_/A _13244_/X _13256_/C VGND VGND VPWR VPWR _13256_/X sky130_fd_sc_hd__and3_4
X_12207_ _12207_/A VGND VGND VPWR VPWR _12207_/Y sky130_fd_sc_hd__inv_2
X_13187_ _13190_/A _18944_/A VGND VGND VPWR VPWR _13188_/C sky130_fd_sc_hd__or2_4
XFILLER_9_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22620__A2 _22422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_72_0_HCLK clkbuf_8_73_0_HCLK/A VGND VGND VPWR VPWR _25113_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16835__B1 _15750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12138_ _24097_/Q _12126_/B _12137_/Y VGND VGND VPWR VPWR _12138_/X sky130_fd_sc_hd__o21a_4
X_19803_ _19802_/Y VGND VGND VPWR VPWR _19803_/X sky130_fd_sc_hd__buf_2
X_17995_ _17995_/A VGND VGND VPWR VPWR _18000_/A sky130_fd_sc_hd__buf_2
XFILLER_111_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22132__A _22132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12069_ _13789_/B _12095_/A VGND VGND VPWR VPWR _16453_/B sky130_fd_sc_hd__or2_4
X_16946_ _16159_/Y _24248_/Q _21426_/A _16927_/X VGND VGND VPWR VPWR _16946_/X sky130_fd_sc_hd__a2bb2o_4
X_19734_ _13288_/B VGND VGND VPWR VPWR _19734_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19665_ _19660_/Y _19663_/X _19664_/X _19663_/X VGND VGND VPWR VPWR _23652_/D sky130_fd_sc_hd__a2bb2o_4
X_16877_ _16875_/Y _16868_/X _16876_/X _16868_/X VGND VGND VPWR VPWR _24396_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18616_ _18616_/A _18616_/B _18616_/C _18615_/X VGND VGND VPWR VPWR _18616_/X sky130_fd_sc_hd__or4_4
X_15828_ _12331_/Y _15826_/X _15756_/X _15826_/X VGND VGND VPWR VPWR _15828_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21690__B _21592_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19596_ _21953_/A _19593_/X _19547_/X _19593_/X VGND VGND VPWR VPWR _19596_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23995__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18547_ _18464_/D _18523_/B _18498_/X _18545_/B VGND VGND VPWR VPWR _18548_/A sky130_fd_sc_hd__a211o_4
X_15759_ _15763_/A VGND VGND VPWR VPWR _15759_/X sky130_fd_sc_hd__buf_2
XFILLER_52_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17012__B1 _24704_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23924__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18478_ _18466_/X _18478_/B VGND VGND VPWR VPWR _18478_/X sky130_fd_sc_hd__or2_4
XANTENNA__25148__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17429_ _24316_/Q VGND VGND VPWR VPWR _17429_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20440_ _20439_/X VGND VGND VPWR VPWR _20443_/B sky130_fd_sc_hd__buf_2
XFILLER_119_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15326__B1 _15318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21211__A _22790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20371_ _21800_/B _20366_/X _11948_/A _20366_/X VGND VGND VPWR VPWR _23391_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12833__A _25361_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22110_ _21306_/A _22106_/X _22109_/X VGND VGND VPWR VPWR _22110_/Y sky130_fd_sc_hd__o21ai_4
X_23090_ _16105_/Y _22551_/X _22843_/X _11766_/Y _22846_/X VGND VGND VPWR VPWR _23090_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__24783__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22041_ _14725_/Y _23671_/Q _14734_/Y _19598_/A VGND VGND VPWR VPWR _22041_/X sky130_fd_sc_hd__o22a_4
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24712__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16826__B1 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16040__A _16060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23992_ _24070_/CLK _20673_/X HRESETn VGND VGND VPWR VPWR _20476_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_56_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22943_ _12849_/D _21438_/X _16941_/Y _22821_/X VGND VGND VPWR VPWR _22943_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19240__B2 _19221_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22874_ _22783_/X _22872_/X _22786_/X _22873_/X VGND VGND VPWR VPWR _22875_/B sky130_fd_sc_hd__o22a_4
XFILLER_43_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23324__B1 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24613_ _24889_/CLK _24613_/D HRESETn VGND VGND VPWR VPWR _22703_/A sky130_fd_sc_hd__dfrtp_4
X_21825_ _21824_/Y _21306_/X _24470_/Q _22873_/B VGND VGND VPWR VPWR _21825_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21756_ _21608_/A _21756_/B VGND VGND VPWR VPWR _21757_/C sky130_fd_sc_hd__or2_4
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24544_ _24561_/CLK _16514_/X HRESETn VGND VGND VPWR VPWR _24544_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25500__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20707_ _13129_/A _13129_/B VGND VGND VPWR VPWR _20707_/X sky130_fd_sc_hd__or2_4
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21687_ _18272_/A _21685_/X _21502_/X _21686_/Y VGND VGND VPWR VPWR _21687_/X sky130_fd_sc_hd__a211o_4
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24475_ _24581_/CLK _24475_/D HRESETn VGND VGND VPWR VPWR _16697_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20638_ _20638_/A _20638_/B VGND VGND VPWR VPWR _20638_/Y sky130_fd_sc_hd__nand2_4
XFILLER_71_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23426_ _23394_/CLK _23426_/D VGND VGND VPWR VPWR _23426_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23357_ _23344_/X VGND VGND VPWR VPWR IRQ[3] sky130_fd_sc_hd__buf_2
X_20569_ _20569_/A VGND VGND VPWR VPWR _20569_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13110_ _13110_/A _13110_/B _13115_/C VGND VGND VPWR VPWR _13110_/X sky130_fd_sc_hd__and3_4
X_22308_ _22308_/A VGND VGND VPWR VPWR _22308_/Y sky130_fd_sc_hd__inv_2
X_14090_ _14089_/X _14026_/Y _14069_/X _13985_/B _14084_/X VGND VGND VPWR VPWR _25215_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_124_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23288_ _23124_/A _23288_/B VGND VGND VPWR VPWR _23288_/Y sky130_fd_sc_hd__nor2_4
XFILLER_69_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13041_ _13041_/A VGND VGND VPWR VPWR _25344_/D sky130_fd_sc_hd__inv_2
X_22239_ _21668_/A _22237_/X _22238_/X VGND VGND VPWR VPWR _22239_/X sky130_fd_sc_hd__and3_4
XANTENNA__14540__A1 scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25027_ _25010_/CLK _15057_/Y HRESETn VGND VGND VPWR VPWR pwm_S6 sky130_fd_sc_hd__dfrtp_4
XANTENNA__23260__C1 _23259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24453__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16817__B1 HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_59_0_HCLK clkbuf_7_58_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16800_ _16799_/Y _16797_/X _15714_/X _16797_/X VGND VGND VPWR VPWR _16800_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17780_ _17805_/A VGND VGND VPWR VPWR _17780_/X sky130_fd_sc_hd__buf_2
X_14992_ _15283_/A _24434_/Q _25000_/Q _14991_/Y VGND VGND VPWR VPWR _14992_/X sky130_fd_sc_hd__a2bb2o_4
X_16731_ _16727_/Y _16730_/X _16376_/X _16730_/X VGND VGND VPWR VPWR _16731_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13943_ _13953_/A _13941_/Y _24954_/Q _13951_/A VGND VGND VPWR VPWR _13943_/X sky130_fd_sc_hd__or4_4
XFILLER_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19450_ _19449_/Y _19447_/X _19404_/X _19447_/X VGND VGND VPWR VPWR _19450_/X sky130_fd_sc_hd__a2bb2o_4
X_16662_ _24489_/Q VGND VGND VPWR VPWR _16662_/Y sky130_fd_sc_hd__inv_2
X_13874_ _21829_/A _13861_/X _21716_/A _13863_/X VGND VGND VPWR VPWR _13874_/X sky130_fd_sc_hd__o22a_4
XFILLER_47_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18401_ _24172_/Q VGND VGND VPWR VPWR _18503_/A sky130_fd_sc_hd__inv_2
XANTENNA__20392__A3 _11862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18990__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23315__B1 _12859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15613_ _22559_/A _15612_/X _11822_/X _15612_/X VGND VGND VPWR VPWR _15613_/X sky130_fd_sc_hd__a2bb2o_4
X_12825_ _25375_/Q VGND VGND VPWR VPWR _12849_/D sky130_fd_sc_hd__inv_2
X_19381_ _17969_/B VGND VGND VPWR VPWR _19381_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20129__B1 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16593_ _16592_/Y _16588_/X _16238_/X _16588_/X VGND VGND VPWR VPWR _16593_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12918__A _12936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18332_ _19219_/C _17486_/X _18331_/X _17451_/Y VGND VGND VPWR VPWR _18332_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11822__A _11821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15544_ _21582_/B VGND VGND VPWR VPWR _15544_/X sky130_fd_sc_hd__buf_2
XFILLER_15_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12756_ _25381_/Q VGND VGND VPWR VPWR _12854_/A sky130_fd_sc_hd__inv_2
XANTENNA__25241__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _24936_/Q VGND VGND VPWR VPWR _11707_/Y sky130_fd_sc_hd__inv_2
X_18263_ _18259_/Y _18262_/Y _16782_/X _18262_/Y VGND VGND VPWR VPWR _18263_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _15473_/Y _15468_/X _15474_/X _15468_/X VGND VGND VPWR VPWR _24941_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12687_ _12674_/X VGND VGND VPWR VPWR _12688_/B sky130_fd_sc_hd__inv_2
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ _16320_/Y _22815_/A _22971_/A _17252_/C VGND VGND VPWR VPWR _17214_/X sky130_fd_sc_hd__a2bb2o_4
X_14426_ _14408_/Y VGND VGND VPWR VPWR _14426_/X sky130_fd_sc_hd__buf_2
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18194_ _15694_/X _18178_/X _18193_/X _24231_/Q _18019_/A VGND VGND VPWR VPWR _18194_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__22127__A _21287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17145_ _17143_/A _17132_/X _17145_/C VGND VGND VPWR VPWR _17145_/X sky130_fd_sc_hd__and3_4
X_14357_ MSO_S3 _14356_/X _25147_/Q _14351_/X VGND VGND VPWR VPWR _14357_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__12653__A _12631_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13308_ _13270_/A _13308_/B VGND VGND VPWR VPWR _13308_/X sky130_fd_sc_hd__or2_4
X_17076_ _17076_/A VGND VGND VPWR VPWR _17076_/Y sky130_fd_sc_hd__inv_2
X_14288_ _25167_/Q VGND VGND VPWR VPWR _14296_/A sky130_fd_sc_hd__inv_2
XANTENNA__16239__A1_N _16237_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16027_ _16002_/X VGND VGND VPWR VPWR _16027_/X sky130_fd_sc_hd__buf_2
XANTENNA__12568__A1_N _12567_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15964__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13239_ _13234_/A VGND VGND VPWR VPWR _13387_/A sky130_fd_sc_hd__buf_2
XFILLER_48_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24194__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16808__B1 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24123__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23003__C1 _23002_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17978_ _18137_/A _17978_/B _17978_/C VGND VGND VPWR VPWR _17979_/C sky130_fd_sc_hd__and3_4
XANTENNA__22797__A _22923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16929_ _21426_/A _16927_/X _22144_/A _16928_/Y VGND VGND VPWR VPWR _16932_/B sky130_fd_sc_hd__a2bb2o_4
X_19717_ _19717_/A VGND VGND VPWR VPWR _19717_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16795__A _16795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19648_ _23657_/Q VGND VGND VPWR VPWR _19648_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25329__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18981__B1 _18961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19579_ _21176_/B _19574_/X _19488_/X _19574_/A VGND VGND VPWR VPWR _23677_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12828__A _25358_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21610_ _14752_/A _18913_/Y VGND VGND VPWR VPWR _21610_/X sky130_fd_sc_hd__or2_4
XFILLER_81_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11732__A _11732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21868__B1 _11844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22590_ _24746_/Q _22590_/B VGND VGND VPWR VPWR _22590_/X sky130_fd_sc_hd__or2_4
XANTENNA__17536__B2 _17565_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21541_ _21333_/A VGND VGND VPWR VPWR _22111_/B sky130_fd_sc_hd__buf_2
XFILLER_138_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24260_ _24682_/CLK _24260_/D HRESETn VGND VGND VPWR VPWR _17754_/A sky130_fd_sc_hd__dfrtp_4
X_21472_ _21477_/A _20375_/Y VGND VGND VPWR VPWR _21472_/X sky130_fd_sc_hd__or2_4
XFILLER_119_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24964__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23211_ _23095_/X _23210_/X _23141_/X _12364_/A _23097_/X VGND VGND VPWR VPWR _23212_/B
+ sky130_fd_sc_hd__a32o_4
X_20423_ _14386_/A _23920_/D _20422_/Y VGND VGND VPWR VPWR _20423_/X sky130_fd_sc_hd__o21a_4
X_24191_ _23377_/CLK _24191_/D HRESETn VGND VGND VPWR VPWR _24191_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12563__A _24847_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16035__A _16060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23142_ _23095_/X _23140_/X _23141_/X _24833_/Q _23097_/X VGND VGND VPWR VPWR _23143_/B
+ sky130_fd_sc_hd__a32o_4
X_20354_ _20354_/A VGND VGND VPWR VPWR _21462_/B sky130_fd_sc_hd__inv_2
X_23073_ _23073_/A _22810_/X _22812_/C VGND VGND VPWR VPWR _23073_/X sky130_fd_sc_hd__and3_4
X_20285_ _20285_/A VGND VGND VPWR VPWR _21915_/B sky130_fd_sc_hd__inv_2
XFILLER_103_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17792__C _17792_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22024_ _22024_/A _19617_/Y VGND VGND VPWR VPWR _22025_/C sky130_fd_sc_hd__or2_4
XANTENNA__22596__B2 _22922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22500__A _22671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23975_ _23978_/CLK _20637_/Y HRESETn VGND VGND VPWR VPWR _20633_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22926_ _16452_/A _22926_/B _22926_/C VGND VGND VPWR VPWR _22926_/X sky130_fd_sc_hd__and3_4
XFILLER_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22857_ _22857_/A _22472_/B VGND VGND VPWR VPWR _22857_/X sky130_fd_sc_hd__or2_4
X_12610_ _12681_/A _12683_/A _12609_/X VGND VGND VPWR VPWR _12666_/A sky130_fd_sc_hd__or3_4
XFILLER_43_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21808_ _21484_/A _21808_/B VGND VGND VPWR VPWR _21808_/X sky130_fd_sc_hd__or2_4
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ _13590_/A _14555_/B VGND VGND VPWR VPWR _14620_/B sky130_fd_sc_hd__and2_4
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22788_ _22783_/X _22785_/X _22786_/X _22787_/X VGND VGND VPWR VPWR _22789_/B sky130_fd_sc_hd__o22a_4
XANTENNA__23331__A _22795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12541_ _25395_/Q VGND VGND VPWR VPWR _12706_/A sky130_fd_sc_hd__inv_2
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24527_ _24557_/CLK _24527_/D HRESETn VGND VGND VPWR VPWR _16560_/A sky130_fd_sc_hd__dfrtp_4
X_21739_ _21739_/A _21019_/A VGND VGND VPWR VPWR _21739_/X sky130_fd_sc_hd__and2_4
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15260_ _15262_/B VGND VGND VPWR VPWR _15261_/B sky130_fd_sc_hd__inv_2
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12472_ _12220_/X _12203_/X _12282_/C _12471_/X VGND VGND VPWR VPWR _12475_/B sky130_fd_sc_hd__or4_4
X_24458_ _25020_/CLK _16742_/X HRESETn VGND VGND VPWR VPWR _24458_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12367__A2_N _24833_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14211_ _14209_/Y _14210_/X _13803_/X _14201_/X VGND VGND VPWR VPWR _14211_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18488__C1 _18487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_22_0_HCLK clkbuf_5_22_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_23409_ _24209_/CLK _20324_/X VGND VGND VPWR VPWR _21978_/C sky130_fd_sc_hd__dfxtp_4
X_15191_ _15191_/A VGND VGND VPWR VPWR _15191_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24389_ _24391_/CLK _17064_/X HRESETn VGND VGND VPWR VPWR _16981_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24634__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ _14102_/A _14102_/B _14102_/A _14102_/B VGND VGND VPWR VPWR _14142_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15784__A _15642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14073_ _14081_/A _14073_/B VGND VGND VPWR VPWR _14073_/X sky130_fd_sc_hd__and2_4
X_18950_ _18949_/Y _18947_/X _17421_/X _18947_/X VGND VGND VPWR VPWR _18950_/X sky130_fd_sc_hd__a2bb2o_4
X_13024_ _13038_/A _13024_/B _13024_/C VGND VGND VPWR VPWR _13024_/X sky130_fd_sc_hd__and3_4
X_17901_ _17889_/X _17898_/Y _17897_/X _17900_/X VGND VGND VPWR VPWR _17901_/X sky130_fd_sc_hd__o22a_4
X_18881_ _23943_/Q _18880_/X VGND VGND VPWR VPWR _18881_/X sky130_fd_sc_hd__or2_4
XFILLER_80_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17832_ _17754_/A _17831_/Y VGND VGND VPWR VPWR _17832_/X sky130_fd_sc_hd__or2_4
XANTENNA__11817__A HWDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17763_ _17786_/A _17762_/X VGND VGND VPWR VPWR _17771_/A sky130_fd_sc_hd__or2_4
X_14975_ _14975_/A VGND VGND VPWR VPWR _14975_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_146_0_HCLK clkbuf_7_73_0_HCLK/X VGND VGND VPWR VPWR _24208_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__25493__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16714_ _16714_/A VGND VGND VPWR VPWR _21582_/A sky130_fd_sc_hd__inv_2
X_19502_ _19502_/A VGND VGND VPWR VPWR _19502_/Y sky130_fd_sc_hd__inv_2
X_13926_ _24961_/Q _13924_/X _13926_/C _13956_/A VGND VGND VPWR VPWR _13942_/C sky130_fd_sc_hd__or4_4
X_17694_ _17689_/X _17694_/B _17681_/X VGND VGND VPWR VPWR _17694_/X sky130_fd_sc_hd__and3_4
XFILLER_48_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25422__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19433_ _18071_/B VGND VGND VPWR VPWR _19433_/Y sky130_fd_sc_hd__inv_2
X_16645_ _16645_/A VGND VGND VPWR VPWR _16658_/A sky130_fd_sc_hd__buf_2
XANTENNA__21026__A _24772_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13857_ _13855_/X _13856_/Y _20466_/B VGND VGND VPWR VPWR _13857_/X sky130_fd_sc_hd__a21o_4
XFILLER_63_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12808_ _12896_/A VGND VGND VPWR VPWR _12887_/A sky130_fd_sc_hd__inv_2
X_19364_ _16781_/X VGND VGND VPWR VPWR _19364_/X sky130_fd_sc_hd__buf_2
XFILLER_76_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16576_ _16574_/Y _16570_/X _16405_/X _16575_/X VGND VGND VPWR VPWR _24521_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13470__C _15652_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13788_ _11723_/Y VGND VGND VPWR VPWR _13789_/D sky130_fd_sc_hd__buf_2
XANTENNA__18715__B1 _18707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18315_ _18295_/A _18314_/Y _18295_/Y _18314_/A VGND VGND VPWR VPWR _18315_/X sky130_fd_sc_hd__o22a_4
X_15527_ _15526_/Y _15524_/X HADDR[8] _15524_/X VGND VGND VPWR VPWR _24920_/D sky130_fd_sc_hd__a2bb2o_4
X_12739_ _12739_/A VGND VGND VPWR VPWR _12739_/Y sky130_fd_sc_hd__inv_2
X_19295_ _19287_/Y VGND VGND VPWR VPWR _19295_/X sky130_fd_sc_hd__buf_2
XANTENNA__15959__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21865__A3 _23005_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18246_ _11686_/Y _18242_/X _16604_/X _18242_/X VGND VGND VPWR VPWR _24221_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15458_ _14280_/X _14251_/A _15446_/A _13897_/X _15452_/X VGND VGND VPWR VPWR _24948_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_129_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_8_0_HCLK_A clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14409_ _14408_/Y VGND VGND VPWR VPWR _14409_/X sky130_fd_sc_hd__buf_2
XANTENNA__22275__B1 _22270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18177_ _18177_/A _18173_/X _18177_/C VGND VGND VPWR VPWR _18178_/C sky130_fd_sc_hd__or3_4
X_15389_ _15389_/A _15388_/X VGND VGND VPWR VPWR _15409_/A sky130_fd_sc_hd__or2_4
XANTENNA__12383__A _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19140__B1 _19071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24375__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17128_ _17156_/A _16985_/Y _16993_/Y _17161_/A VGND VGND VPWR VPWR _17128_/X sky130_fd_sc_hd__or4_4
XFILLER_117_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24304__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17059_ _17050_/A _17050_/D VGND VGND VPWR VPWR _17060_/B sky130_fd_sc_hd__or2_4
X_20070_ _20064_/X _18326_/X _15836_/X _13312_/B _20066_/X VGND VGND VPWR VPWR _23505_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_42_0_HCLK clkbuf_7_42_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_42_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17414__A _21355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20972_ _24108_/Q _24106_/Q VGND VGND VPWR VPWR _20972_/X sky130_fd_sc_hd__and2_4
X_23760_ _23828_/CLK _19344_/X VGND VGND VPWR VPWR _18118_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__25163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22711_ _22711_/A _22711_/B _22705_/X _22710_/X VGND VGND VPWR VPWR _22711_/X sky130_fd_sc_hd__or4_4
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23691_ _23384_/CLK _19542_/X VGND VGND VPWR VPWR _23691_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25430_ _25425_/CLK _25430_/D HRESETn VGND VGND VPWR VPWR _25430_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_94_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22642_ _22642_/A VGND VGND VPWR VPWR _22642_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14440__B1 _14414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12277__B _12277_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22502__B2 _22790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23151__A _22654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25361_ _25330_/CLK _25361_/D HRESETn VGND VGND VPWR VPWR _25361_/Q sky130_fd_sc_hd__dfrtp_4
X_22573_ _24412_/Q _22523_/X _22524_/X _22572_/X VGND VGND VPWR VPWR _22574_/C sky130_fd_sc_hd__a211o_4
XFILLER_22_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24312_ _24885_/CLK _17444_/X HRESETn VGND VGND VPWR VPWR _24312_/Q sky130_fd_sc_hd__dfrtp_4
X_21524_ _22489_/A VGND VGND VPWR VPWR _21524_/X sky130_fd_sc_hd__buf_2
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25292_ _25478_/CLK _25292_/D HRESETn VGND VGND VPWR VPWR SCLK_S2 sky130_fd_sc_hd__dfstp_4
XFILLER_72_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21455_ _21455_/A VGND VGND VPWR VPWR _21456_/A sky130_fd_sc_hd__buf_2
X_24243_ _24288_/CLK _24243_/D HRESETn VGND VGND VPWR VPWR _24243_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19131__B1 _19018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20406_ _20404_/Y _20400_/X _11842_/A _20405_/X VGND VGND VPWR VPWR _23376_/D sky130_fd_sc_hd__a2bb2o_4
X_24174_ _24171_/CLK _24174_/D HRESETn VGND VGND VPWR VPWR _18414_/A sky130_fd_sc_hd__dfrtp_4
X_21386_ _21391_/A _21384_/X _21386_/C VGND VGND VPWR VPWR _21386_/X sky130_fd_sc_hd__and3_4
XANTENNA__24045__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20337_ _20337_/A VGND VGND VPWR VPWR _22332_/B sky130_fd_sc_hd__inv_2
XANTENNA__19076__A _19062_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23125_ _22795_/A VGND VGND VPWR VPWR _23208_/A sky130_fd_sc_hd__buf_2
X_23056_ _23056_/A _23055_/X VGND VGND VPWR VPWR _23066_/B sky130_fd_sc_hd__nor2_4
X_20268_ _20268_/A VGND VGND VPWR VPWR _20268_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23230__A2 _22988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22007_ _22025_/A _22007_/B _22006_/X VGND VGND VPWR VPWR _22007_/X sky130_fd_sc_hd__and3_4
XFILLER_89_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20199_ _21882_/B _20196_/X _19787_/A _20196_/X VGND VGND VPWR VPWR _20199_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13852__A _23989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_219_0_HCLK clkbuf_8_219_0_HCLK/A VGND VGND VPWR VPWR _24447_/CLK sky130_fd_sc_hd__clkbuf_1
X_14760_ _13744_/A VGND VGND VPWR VPWR _14770_/B sky130_fd_sc_hd__buf_2
X_11972_ _11647_/X _11650_/A VGND VGND VPWR VPWR _11972_/X sky130_fd_sc_hd__or2_4
X_23958_ _23989_/CLK _20473_/X HRESETn VGND VGND VPWR VPWR _21351_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22741__A1 _22476_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13711_ _13691_/B _13707_/X _13710_/Y _13703_/X _25278_/Q VGND VGND VPWR VPWR _13711_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22741__B2 _22480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22909_ _22764_/A VGND VGND VPWR VPWR _22909_/X sky130_fd_sc_hd__buf_2
X_14691_ _14691_/A VGND VGND VPWR VPWR _21391_/A sky130_fd_sc_hd__buf_2
X_23889_ _23854_/CLK _23889_/D VGND VGND VPWR VPWR _23889_/Q sky130_fd_sc_hd__dfxtp_4
X_16430_ _15112_/Y _16426_/X _16143_/X _16429_/X VGND VGND VPWR VPWR _16430_/X sky130_fd_sc_hd__a2bb2o_4
X_13642_ _13640_/X _13642_/B VGND VGND VPWR VPWR _13642_/X sky130_fd_sc_hd__or2_4
XFILLER_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23297__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24886__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16361_ _21531_/A VGND VGND VPWR VPWR _16361_/Y sky130_fd_sc_hd__inv_2
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _13573_/A VGND VGND VPWR VPWR _13573_/Y sky130_fd_sc_hd__inv_2
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14982__B2 _16850_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18100_ _18196_/A _23752_/Q VGND VGND VPWR VPWR _18102_/B sky130_fd_sc_hd__or2_4
XANTENNA__24815__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15312_ _24994_/Q _15312_/B VGND VGND VPWR VPWR _15314_/B sky130_fd_sc_hd__or2_4
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _12524_/A VGND VGND VPWR VPWR _12524_/Y sky130_fd_sc_hd__inv_2
X_19080_ _19079_/Y _19076_/X _19056_/X _19076_/X VGND VGND VPWR VPWR _19080_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _16291_/Y _16289_/X _15942_/X _16289_/X VGND VGND VPWR VPWR _16292_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12915__B _12903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18031_ _18137_/A _18031_/B _18031_/C VGND VGND VPWR VPWR _18032_/C sky130_fd_sc_hd__and3_4
X_15243_ _15216_/A _15243_/B _15242_/X VGND VGND VPWR VPWR _25008_/D sky130_fd_sc_hd__and3_4
X_12455_ _12249_/X _12455_/B VGND VGND VPWR VPWR _12456_/C sky130_fd_sc_hd__or2_4
XFILLER_138_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15174_ _15199_/A VGND VGND VPWR VPWR _15174_/X sky130_fd_sc_hd__buf_2
XFILLER_67_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12386_ _12385_/X VGND VGND VPWR VPWR _12387_/B sky130_fd_sc_hd__inv_2
X_14125_ _14125_/A VGND VGND VPWR VPWR _14125_/X sky130_fd_sc_hd__buf_2
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19982_ _19991_/A VGND VGND VPWR VPWR _19982_/X sky130_fd_sc_hd__buf_2
XANTENNA__12931__A _12602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16403__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22124__B _22836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14056_ _14056_/A VGND VGND VPWR VPWR _14078_/A sky130_fd_sc_hd__buf_2
X_18933_ _18932_/Y _18930_/X _16782_/X _18930_/X VGND VGND VPWR VPWR _23905_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13007_ _13026_/A VGND VGND VPWR VPWR _13010_/A sky130_fd_sc_hd__buf_2
XFILLER_79_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_29_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_58_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18864_ _18860_/X _18861_/X _18864_/C _18864_/D VGND VGND VPWR VPWR _18865_/D sky130_fd_sc_hd__or4_4
XFILLER_79_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17815_ _17834_/A _17815_/B _17815_/C VGND VGND VPWR VPWR _17815_/X sky130_fd_sc_hd__and3_4
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18795_ _18792_/B _18792_/C VGND VGND VPWR VPWR _18796_/A sky130_fd_sc_hd__or2_4
XANTENNA__15998__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19189__B1 _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19472__A2_N _19471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17746_ _21048_/A VGND VGND VPWR VPWR _17747_/D sky130_fd_sc_hd__inv_2
X_14958_ _15227_/A VGND VGND VPWR VPWR _15219_/B sky130_fd_sc_hd__inv_2
XFILLER_54_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13909_ _13909_/A _24952_/Q _13909_/C _24950_/Q VGND VGND VPWR VPWR _13909_/X sky130_fd_sc_hd__or4_4
XFILLER_130_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17677_ _17652_/X _17674_/B _17677_/C VGND VGND VPWR VPWR _17677_/X sky130_fd_sc_hd__and3_4
X_14889_ _14888_/Y _24432_/Q _14888_/Y _24432_/Q VGND VGND VPWR VPWR _14889_/X sky130_fd_sc_hd__a2bb2o_4
X_16628_ _16173_/A _14766_/X _16624_/X _13740_/A _16627_/X VGND VGND VPWR VPWR _24501_/D
+ sky130_fd_sc_hd__a32o_4
X_19416_ _19414_/Y _19415_/X _19370_/X _19415_/X VGND VGND VPWR VPWR _19416_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16559_ _16557_/Y _16558_/X _16297_/X _16558_/X VGND VGND VPWR VPWR _16559_/X sky130_fd_sc_hd__a2bb2o_4
X_19347_ _19345_/Y _19346_/X _19212_/X _19346_/X VGND VGND VPWR VPWR _23759_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22496__B1 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24556__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19278_ _19278_/A VGND VGND VPWR VPWR _19278_/X sky130_fd_sc_hd__buf_2
XFILLER_31_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18229_ _17448_/X VGND VGND VPWR VPWR _18230_/B sky130_fd_sc_hd__buf_2
XFILLER_15_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19113__B1 _18997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21240_ _21372_/A VGND VGND VPWR VPWR _21240_/X sky130_fd_sc_hd__buf_2
XFILLER_102_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21171_ _21165_/X _21170_/X _17719_/Y VGND VGND VPWR VPWR _21171_/X sky130_fd_sc_hd__o21a_4
XFILLER_117_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20122_ _23485_/Q VGND VGND VPWR VPWR _20122_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20053_ _21904_/B _20050_/X _19787_/X _20050_/X VGND VGND VPWR VPWR _20053_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24930_ _24930_/CLK _24930_/D HRESETn VGND VGND VPWR VPWR _11727_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25344__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16055__A1_N _16054_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15989__B1 _24735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24861_ _24847_/CLK _24861_/D HRESETn VGND VGND VPWR VPWR _12533_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21592__C _21578_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17144__A _17038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23812_ _23818_/CLK _19199_/X VGND VGND VPWR VPWR _19195_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_27_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24792_ _24792_/CLK _15881_/X HRESETn VGND VGND VPWR VPWR _24792_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13464__B2 _13195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22723__A1 _24448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_192_0_HCLK clkbuf_7_96_0_HCLK/X VGND VGND VPWR VPWR _24334_/CLK sky130_fd_sc_hd__clkbuf_1
X_23743_ _23446_/CLK _19393_/X VGND VGND VPWR VPWR _18133_/B sky130_fd_sc_hd__dfxtp_4
X_20955_ _12006_/A _20955_/B VGND VGND VPWR VPWR _24087_/D sky130_fd_sc_hd__and2_4
XPHY_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_49_0_HCLK clkbuf_8_49_0_HCLK/A VGND VGND VPWR VPWR _25290_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23674_ _23384_/CLK _23674_/D VGND VGND VPWR VPWR _21963_/C sky130_fd_sc_hd__dfxtp_4
X_20886_ _20913_/A VGND VGND VPWR VPWR _20886_/X sky130_fd_sc_hd__buf_2
XPHY_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25413_ _25400_/CLK _12655_/X HRESETn VGND VGND VPWR VPWR _25413_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22625_ _22549_/A _22625_/B VGND VGND VPWR VPWR _22625_/Y sky130_fd_sc_hd__nand2_4
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19352__B1 _19307_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24297__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25344_ _23370_/CLK _25344_/D HRESETn VGND VGND VPWR VPWR _25344_/Q sky130_fd_sc_hd__dfrtp_4
X_22556_ _22556_/A _21085_/A VGND VGND VPWR VPWR _22556_/X sky130_fd_sc_hd__or2_4
XANTENNA__16166__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24226__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16623__A1_N _16622_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21507_ _21160_/X VGND VGND VPWR VPWR _21507_/Y sky130_fd_sc_hd__inv_2
X_25275_ _25279_/CLK _25275_/D HRESETn VGND VGND VPWR VPWR _11667_/A sky130_fd_sc_hd__dfrtp_4
X_22487_ _22475_/X _22482_/Y _22483_/X _22486_/X VGND VGND VPWR VPWR _22487_/X sky130_fd_sc_hd__a2bb2o_4
X_12240_ _12230_/X _12240_/B _12236_/X _12239_/X VGND VGND VPWR VPWR _12272_/A sky130_fd_sc_hd__or4_4
X_24226_ _24346_/CLK _24226_/D HRESETn VGND VGND VPWR VPWR _24226_/Q sky130_fd_sc_hd__dfrtp_4
X_21438_ _21009_/X VGND VGND VPWR VPWR _21438_/X sky130_fd_sc_hd__buf_2
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22225__A _21192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12171_ _25453_/Q VGND VGND VPWR VPWR SSn_S3 sky130_fd_sc_hd__inv_2
X_21369_ _18230_/A _21367_/X _13782_/X _21368_/X VGND VGND VPWR VPWR _21369_/X sky130_fd_sc_hd__a211o_4
X_24157_ _24159_/CLK _24157_/D HRESETn VGND VGND VPWR VPWR _24157_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23108_ _23106_/X _23107_/X _23040_/X _16012_/A _22972_/X VGND VGND VPWR VPWR _23108_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17038__B _17038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24088_ _25301_/CLK _20956_/X HRESETn VGND VGND VPWR VPWR _24088_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15930_ _15795_/A VGND VGND VPWR VPWR _15930_/X sky130_fd_sc_hd__buf_2
XANTENNA__22411__B1 _12542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23039_ _23039_/A _22898_/X VGND VGND VPWR VPWR _23039_/X sky130_fd_sc_hd__or2_4
XANTENNA__21537__A2_N _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25085__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15861_ _21026_/B VGND VGND VPWR VPWR _15931_/B sky130_fd_sc_hd__buf_2
XFILLER_27_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25014__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17600_ _17560_/Y _17582_/X _17600_/C _17600_/D VGND VGND VPWR VPWR _17600_/X sky130_fd_sc_hd__or4_4
X_14812_ _14803_/C VGND VGND VPWR VPWR _14819_/A sky130_fd_sc_hd__inv_2
XFILLER_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16641__A1 _15824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18580_ _18580_/A VGND VGND VPWR VPWR _18581_/B sky130_fd_sc_hd__inv_2
X_15792_ _15817_/A VGND VGND VPWR VPWR _15793_/A sky130_fd_sc_hd__buf_2
XFILLER_79_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17531_ _11802_/Y _24292_/Q _11802_/Y _24292_/Q VGND VGND VPWR VPWR _17531_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14743_ _14742_/Y _14723_/Y _22038_/A _14722_/X VGND VGND VPWR VPWR _14743_/X sky130_fd_sc_hd__o22a_4
X_11955_ _19632_/A VGND VGND VPWR VPWR _11955_/X sky130_fd_sc_hd__buf_2
XFILLER_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19591__B1 _19404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18394__B2 _24172_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17462_ _24196_/Q VGND VGND VPWR VPWR _17462_/Y sky130_fd_sc_hd__inv_2
X_14674_ _25057_/Q VGND VGND VPWR VPWR _21781_/A sky130_fd_sc_hd__inv_2
X_11886_ _11886_/A VGND VGND VPWR VPWR _11886_/Y sky130_fd_sc_hd__inv_2
X_16413_ _16381_/A VGND VGND VPWR VPWR _16433_/A sky130_fd_sc_hd__buf_2
X_19201_ _19200_/Y _19198_/X _19133_/X _19198_/X VGND VGND VPWR VPWR _23811_/D sky130_fd_sc_hd__a2bb2o_4
X_13625_ _14658_/A VGND VGND VPWR VPWR _19152_/D sky130_fd_sc_hd__buf_2
XFILLER_73_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17393_ _20633_/A _17392_/X VGND VGND VPWR VPWR _20638_/B sky130_fd_sc_hd__or2_4
XFILLER_20_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19132_ _19132_/A VGND VGND VPWR VPWR _19132_/Y sky130_fd_sc_hd__inv_2
X_16344_ _16342_/Y _16337_/X _16143_/X _16343_/X VGND VGND VPWR VPWR _24608_/D sky130_fd_sc_hd__a2bb2o_4
X_13556_ _22726_/A _25085_/Q _22726_/A _25085_/Q VGND VGND VPWR VPWR _13564_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12507_ _13042_/A VGND VGND VPWR VPWR _13026_/A sky130_fd_sc_hd__inv_2
X_19063_ _19062_/Y VGND VGND VPWR VPWR _19063_/X sky130_fd_sc_hd__buf_2
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16275_ _22884_/B VGND VGND VPWR VPWR _22671_/A sky130_fd_sc_hd__buf_2
X_13487_ _13486_/Y _13482_/X _11853_/X _13482_/X VGND VGND VPWR VPWR _25307_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18014_ _18010_/A VGND VGND VPWR VPWR _18056_/A sky130_fd_sc_hd__buf_2
X_15226_ _15223_/B VGND VGND VPWR VPWR _15227_/B sky130_fd_sc_hd__inv_2
X_12438_ _12433_/A _12433_/B _12402_/X _12434_/Y VGND VGND VPWR VPWR _12438_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22135__A _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15157_ _24991_/Q _15145_/Y _15389_/A _24571_/Q VGND VGND VPWR VPWR _15161_/C sky130_fd_sc_hd__a2bb2o_4
X_12369_ _25342_/Q VGND VGND VPWR VPWR _12990_/B sky130_fd_sc_hd__inv_2
XFILLER_113_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14108_ _14108_/A VGND VGND VPWR VPWR _14108_/X sky130_fd_sc_hd__buf_2
XFILLER_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15088_ _24973_/Q _15086_/Y _15087_/Y _24593_/Q VGND VGND VPWR VPWR _15088_/X sky130_fd_sc_hd__a2bb2o_4
X_19965_ _19963_/Y _19964_/X _19629_/X _19964_/X VGND VGND VPWR VPWR _19965_/X sky130_fd_sc_hd__a2bb2o_4
X_14039_ _13975_/A _14007_/X VGND VGND VPWR VPWR _14039_/Y sky130_fd_sc_hd__nand2_4
X_18916_ _18916_/A VGND VGND VPWR VPWR _21384_/B sky130_fd_sc_hd__inv_2
X_19896_ _19894_/Y _19890_/X _19618_/X _19895_/X VGND VGND VPWR VPWR _23570_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18847_ _21837_/A _18678_/Y _24540_/Q _18782_/X VGND VGND VPWR VPWR _18849_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25154__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18778_ _18692_/B _18773_/B _18733_/X _18774_/Y VGND VGND VPWR VPWR _18778_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_202_0_HCLK clkbuf_8_203_0_HCLK/A VGND VGND VPWR VPWR _25354_/CLK sky130_fd_sc_hd__clkbuf_1
X_17729_ _17729_/A VGND VGND VPWR VPWR _17729_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24737__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_8_0_HCLK clkbuf_7_4_0_HCLK/X VGND VGND VPWR VPWR _23498_/CLK sky130_fd_sc_hd__clkbuf_1
X_20740_ _20740_/A _20740_/B VGND VGND VPWR VPWR _20740_/X sky130_fd_sc_hd__or2_4
XFILLER_90_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21214__A _16719_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20671_ _20481_/X _20488_/X _20602_/X VGND VGND VPWR VPWR _20671_/X sky130_fd_sc_hd__o21a_4
XFILLER_91_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11740__A _11739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24390__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22410_ _24779_/Q _21073_/B VGND VGND VPWR VPWR _22410_/X sky130_fd_sc_hd__or2_4
XANTENNA__16148__B1 _16147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21141__B1 _14881_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23390_ _23533_/CLK _23390_/D VGND VGND VPWR VPWR _23390_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22341_ _21917_/X _22341_/B _22340_/X VGND VGND VPWR VPWR _22341_/X sky130_fd_sc_hd__and3_4
XANTENNA__21692__A1 _21512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21692__B2 _21428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22272_ _21530_/X VGND VGND VPWR VPWR _22272_/X sky130_fd_sc_hd__buf_2
XFILLER_136_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25060_ _25044_/CLK _14668_/X HRESETn VGND VGND VPWR VPWR _13624_/A sky130_fd_sc_hd__dfrtp_4
X_21223_ _21252_/A _21223_/B VGND VGND VPWR VPWR _21226_/B sky130_fd_sc_hd__or2_4
X_24011_ _24909_/CLK _20742_/X HRESETn VGND VGND VPWR VPWR _20740_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25525__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21154_ _16855_/Y _21154_/B VGND VGND VPWR VPWR _21157_/B sky130_fd_sc_hd__or2_4
XFILLER_137_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20105_ _20105_/A VGND VGND VPWR VPWR _20105_/X sky130_fd_sc_hd__buf_2
XFILLER_132_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22699__B _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21085_ _21085_/A VGND VGND VPWR VPWR _22587_/B sky130_fd_sc_hd__buf_2
XFILLER_59_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14882__B1 _14881_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22944__A1 _12433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20036_ _20036_/A VGND VGND VPWR VPWR _20036_/X sky130_fd_sc_hd__buf_2
X_24913_ _24923_/CLK _15541_/X HRESETn VGND VGND VPWR VPWR _24913_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_12_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_86_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16623__B2 _16545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24844_ _24847_/CLK _24844_/D HRESETn VGND VGND VPWR VPWR _12552_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_37_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21108__B _21108_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24775_ _24811_/CLK _15907_/X HRESETn VGND VGND VPWR VPWR _24775_/Q sky130_fd_sc_hd__dfrtp_4
X_21987_ _17909_/A _20335_/Y _21987_/C VGND VGND VPWR VPWR _21987_/X sky130_fd_sc_hd__and3_4
XFILLER_54_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24478__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11739_/X VGND VGND VPWR VPWR _11750_/A sky130_fd_sc_hd__buf_2
XPHY_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23726_ _23722_/CLK _23726_/D VGND VGND VPWR VPWR _18172_/B sky130_fd_sc_hd__dfxtp_4
X_20938_ _24057_/Q VGND VGND VPWR VPWR _20939_/A sky130_fd_sc_hd__inv_2
XANTENNA__16387__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23323__B _22832_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24407__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _24224_/Q VGND VGND VPWR VPWR _11671_/Y sky130_fd_sc_hd__inv_2
XPHY_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23657_ _24197_/CLK _19649_/X VGND VGND VPWR VPWR _23657_/Q sky130_fd_sc_hd__dfxtp_4
X_20869_ _20860_/X _20868_/X _24477_/Q _20865_/X VGND VGND VPWR VPWR _24040_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12261__A1_N _12252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13156_/X _13410_/B _13409_/X VGND VGND VPWR VPWR _13410_/X sky130_fd_sc_hd__and3_4
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16139__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22608_ _22608_/A _22522_/B VGND VGND VPWR VPWR _22608_/X sky130_fd_sc_hd__or2_4
X_14390_ _20420_/B VGND VGND VPWR VPWR _20496_/D sky130_fd_sc_hd__inv_2
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23588_ _23498_/CLK _23588_/D VGND VGND VPWR VPWR _23588_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24060__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13341_ _13373_/A _13341_/B VGND VGND VPWR VPWR _13341_/X sky130_fd_sc_hd__or2_4
XFILLER_128_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21683__A1 _20331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25327_ _24836_/CLK _25327_/D HRESETn VGND VGND VPWR VPWR _13102_/A sky130_fd_sc_hd__dfrtp_4
X_22539_ _22539_/A _16373_/A VGND VGND VPWR VPWR _22539_/X sky130_fd_sc_hd__or2_4
XANTENNA__22880__B1 _22798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21683__B2 _22390_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16060_ _16060_/A VGND VGND VPWR VPWR _16060_/X sky130_fd_sc_hd__buf_2
X_13272_ _13310_/A _13272_/B VGND VGND VPWR VPWR _13272_/X sky130_fd_sc_hd__or2_4
X_25258_ _25070_/CLK _25258_/D HRESETn VGND VGND VPWR VPWR _25258_/Q sky130_fd_sc_hd__dfrtp_4
X_15011_ _24997_/Q _24435_/Q _15278_/A _15010_/Y VGND VGND VPWR VPWR _15012_/D sky130_fd_sc_hd__o22a_4
X_12223_ _25422_/Q VGND VGND VPWR VPWR _12499_/A sky130_fd_sc_hd__inv_2
XANTENNA__21435__A1 _21280_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24209_ _24209_/CLK _18268_/X HRESETn VGND VGND VPWR VPWR _24209_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21435__B2 _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25266__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25189_ _25192_/CLK _14217_/X HRESETn VGND VGND VPWR VPWR _20664_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_118_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12154_ _12152_/A _12153_/A _12152_/Y _12153_/Y VGND VGND VPWR VPWR _12154_/X sky130_fd_sc_hd__o22a_4
XFILLER_29_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22392__A1_N _21270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15792__A _15817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19750_ _19728_/A _17472_/A _18922_/X VGND VGND VPWR VPWR _19750_/X sky130_fd_sc_hd__or3_4
X_12085_ _25468_/Q VGND VGND VPWR VPWR _12085_/Y sky130_fd_sc_hd__inv_2
X_16962_ _16012_/Y _24385_/Q _16012_/Y _24385_/Q VGND VGND VPWR VPWR _16962_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22402__B _22266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18701_ _18599_/X _18701_/B VGND VGND VPWR VPWR _18701_/Y sky130_fd_sc_hd__nand2_4
XFILLER_77_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15913_ _14769_/X _15911_/Y _15912_/X VGND VGND VPWR VPWR _15913_/X sky130_fd_sc_hd__o21a_4
X_16893_ _22183_/A _17867_/A _16098_/Y _17785_/A VGND VGND VPWR VPWR _16893_/X sky130_fd_sc_hd__a2bb2o_4
X_19681_ _19680_/Y _19676_/X _19658_/X _19676_/A VGND VGND VPWR VPWR _19681_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19800__B2 _19793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11825__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15844_ _15646_/X _15765_/X _15774_/X _21006_/B _15843_/X VGND VGND VPWR VPWR _15844_/X
+ sky130_fd_sc_hd__a32o_4
X_18632_ _24511_/Q _18630_/A _16599_/Y _18792_/A VGND VGND VPWR VPWR _18632_/X sky130_fd_sc_hd__o22a_4
XFILLER_18_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15968__A3 HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15775_ _15777_/A _15843_/A VGND VGND VPWR VPWR _15775_/X sky130_fd_sc_hd__or2_4
X_18563_ _18411_/Y _18575_/B VGND VGND VPWR VPWR _18576_/B sky130_fd_sc_hd__or2_4
XFILLER_79_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12987_ _25343_/Q VGND VGND VPWR VPWR _13048_/A sky130_fd_sc_hd__inv_2
XFILLER_92_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24830__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14726_ _14725_/Y _14708_/X _25054_/Q _14707_/A VGND VGND VPWR VPWR _14726_/X sky130_fd_sc_hd__o22a_4
X_17514_ _17514_/A _17509_/X _17514_/C _17513_/X VGND VGND VPWR VPWR _17514_/X sky130_fd_sc_hd__or4_4
XFILLER_18_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11938_ _19622_/A VGND VGND VPWR VPWR _11938_/Y sky130_fd_sc_hd__inv_2
X_18494_ _18481_/B _18491_/X VGND VGND VPWR VPWR _18494_/X sky130_fd_sc_hd__or2_4
XFILLER_45_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24148__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17445_ _25539_/Q _17445_/B _17445_/C VGND VGND VPWR VPWR _17474_/A sky130_fd_sc_hd__or3_4
X_14657_ _14656_/Y VGND VGND VPWR VPWR _19038_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_32_0_HCLK clkbuf_7_16_0_HCLK/X VGND VGND VPWR VPWR _23805_/CLK sky130_fd_sc_hd__clkbuf_1
X_11869_ _25505_/Q _11869_/B VGND VGND VPWR VPWR _11869_/X sky130_fd_sc_hd__and2_4
XANTENNA__19316__B1 _19291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_95_0_HCLK clkbuf_8_95_0_HCLK/A VGND VGND VPWR VPWR _24133_/CLK sky130_fd_sc_hd__clkbuf_1
X_13608_ _13626_/B VGND VGND VPWR VPWR _13609_/B sky130_fd_sc_hd__inv_2
X_17376_ _17206_/X _17347_/B VGND VGND VPWR VPWR _17377_/B sky130_fd_sc_hd__or2_4
X_14588_ _14573_/A _14586_/X _14587_/X _13770_/X _25081_/Q VGND VGND VPWR VPWR _14588_/X
+ sky130_fd_sc_hd__a32o_4
X_16327_ _24614_/Q VGND VGND VPWR VPWR _16327_/Y sky130_fd_sc_hd__inv_2
X_19115_ _19114_/Y _19112_/X _19071_/X _19112_/X VGND VGND VPWR VPWR _23841_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_14_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13539_ _24771_/Q VGND VGND VPWR VPWR _15677_/A sky130_fd_sc_hd__inv_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19046_ _19044_/Y _19040_/X _18997_/X _19045_/X VGND VGND VPWR VPWR _19046_/X sky130_fd_sc_hd__a2bb2o_4
X_16258_ _21836_/A VGND VGND VPWR VPWR _16258_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15209_ _15209_/A _15239_/A _15209_/C _15171_/B VGND VGND VPWR VPWR _15210_/C sky130_fd_sc_hd__or4_4
X_16189_ _23291_/A VGND VGND VPWR VPWR _16189_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19948_ _19947_/Y _19943_/X _19885_/X _19943_/A VGND VGND VPWR VPWR _19948_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24989__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19879_ _19879_/A VGND VGND VPWR VPWR _21650_/B sky130_fd_sc_hd__inv_2
XANTENNA__24918__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21910_ _14716_/A _21902_/X _21909_/X VGND VGND VPWR VPWR _21910_/X sky130_fd_sc_hd__or3_4
XANTENNA__11735__A _21314_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22890_ _22868_/X _22871_/X _22875_/Y _22889_/X VGND VGND VPWR VPWR HRDATA[18] sky130_fd_sc_hd__a211o_4
XANTENNA__18651__A1_N _16585_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21841_ _21841_/A _22111_/B VGND VGND VPWR VPWR _21841_/Y sky130_fd_sc_hd__nand2_4
XFILLER_71_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24571__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24560_ _24557_/CLK _16475_/X HRESETn VGND VGND VPWR VPWR _24560_/Q sky130_fd_sc_hd__dfrtp_4
X_21772_ _21596_/A _21772_/B VGND VGND VPWR VPWR _21772_/X sky130_fd_sc_hd__or2_4
XFILLER_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24500__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23511_ _25055_/CLK _23511_/D VGND VGND VPWR VPWR _20056_/A sky130_fd_sc_hd__dfxtp_4
X_20723_ _24007_/Q _13130_/B _20722_/Y VGND VGND VPWR VPWR _20723_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24491_ _24447_/CLK _24491_/D HRESETn VGND VGND VPWR VPWR _24491_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23442_ _23441_/CLK _23442_/D VGND VGND VPWR VPWR _13266_/B sky130_fd_sc_hd__dfxtp_4
X_20654_ _25186_/Q _17404_/A VGND VGND VPWR VPWR _20657_/B sky130_fd_sc_hd__or2_4
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_3_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20585_ _14394_/A _20582_/X _20584_/X VGND VGND VPWR VPWR _23942_/D sky130_fd_sc_hd__and3_4
XANTENNA__19349__A _19055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23373_ _23904_/CLK _23373_/D VGND VGND VPWR VPWR _13376_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_128_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25112_ _25101_/CLK _25112_/D HRESETn VGND VGND VPWR VPWR _25112_/Q sky130_fd_sc_hd__dfrtp_4
X_22324_ _21332_/Y _22309_/X _22311_/X _22315_/Y _22323_/X VGND VGND VPWR VPWR _22383_/C
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__22614__B1 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25043_ _25043_/CLK _14821_/X HRESETn VGND VGND VPWR VPWR _14805_/A sky130_fd_sc_hd__dfrtp_4
X_22255_ _18291_/X _22251_/X _22255_/C VGND VGND VPWR VPWR _22255_/X sky130_fd_sc_hd__or3_4
X_21206_ _21205_/X VGND VGND VPWR VPWR _21207_/C sky130_fd_sc_hd__inv_2
X_22186_ _22186_/A _22186_/B _22186_/C VGND VGND VPWR VPWR _22187_/D sky130_fd_sc_hd__and3_4
XFILLER_117_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18604__A1_N _16560_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21137_ _21133_/X _21137_/B VGND VGND VPWR VPWR _21137_/X sky130_fd_sc_hd__and2_4
XFILLER_78_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23318__B _16795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21068_ _21154_/B VGND VGND VPWR VPWR _21069_/A sky130_fd_sc_hd__buf_2
XFILLER_87_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21119__A _21119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24659__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12910_ _12849_/D _12905_/B _12874_/X _12906_/Y VGND VGND VPWR VPWR _12911_/A sky130_fd_sc_hd__a211o_4
X_20019_ _19885_/A VGND VGND VPWR VPWR _20019_/X sky130_fd_sc_hd__buf_2
XFILLER_111_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13890_ _24961_/Q _13924_/A _13889_/X VGND VGND VPWR VPWR _13958_/D sky130_fd_sc_hd__or3_4
XFILLER_74_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12841_ _12749_/Y _12841_/B VGND VGND VPWR VPWR _12841_/X sky130_fd_sc_hd__or2_4
X_24827_ _24868_/CLK _15811_/X HRESETn VGND VGND VPWR VPWR _24827_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13860__A _23990_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15560_ _15560_/A VGND VGND VPWR VPWR _15580_/A sky130_fd_sc_hd__inv_2
XANTENNA__17332__A _17252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12772_ _12772_/A VGND VGND VPWR VPWR _12772_/Y sky130_fd_sc_hd__inv_2
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24758_ _24821_/CLK _15951_/X HRESETn VGND VGND VPWR VPWR _24758_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24241__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14510_/X VGND VGND VPWR VPWR _14511_/X sky130_fd_sc_hd__buf_2
XPHY_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _24914_/Q VGND VGND VPWR VPWR _11723_/Y sky130_fd_sc_hd__inv_2
XPHY_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23709_ _23396_/CLK _19489_/X VGND VGND VPWR VPWR _23709_/Q sky130_fd_sc_hd__dfxtp_4
X_15491_ _15490_/X VGND VGND VPWR VPWR _15491_/X sky130_fd_sc_hd__buf_2
XPHY_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_19_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24689_ _24689_/CLK _16114_/X HRESETn VGND VGND VPWR VPWR _22976_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17230_/A _17216_/X _17224_/X _17230_/D VGND VGND VPWR VPWR _17231_/B sky130_fd_sc_hd__or4_4
XPHY_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14436_/Y VGND VGND VPWR VPWR _14442_/X sky130_fd_sc_hd__buf_2
XFILLER_80_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11654_/A _11654_/B _11654_/C VGND VGND VPWR VPWR _11655_/A sky130_fd_sc_hd__and3_4
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16780__B1 _16528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17161_ _17161_/A VGND VGND VPWR VPWR _17162_/B sky130_fd_sc_hd__inv_2
XFILLER_31_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14373_ _25140_/Q VGND VGND VPWR VPWR _14373_/Y sky130_fd_sc_hd__inv_2
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20778__A1_N _20770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15002__D _15002_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25447__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16112_ _22976_/A VGND VGND VPWR VPWR _16112_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13324_ _13246_/X _23633_/Q VGND VGND VPWR VPWR _13324_/X sky130_fd_sc_hd__or2_4
XFILLER_70_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17092_ _17034_/X _17091_/X VGND VGND VPWR VPWR _17092_/X sky130_fd_sc_hd__or2_4
XANTENNA__16532__B1 _16355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16043_ _16042_/Y _16040_/X _11809_/X _16040_/X VGND VGND VPWR VPWR _24716_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13255_ _13162_/X _13255_/B _13254_/X VGND VGND VPWR VPWR _13256_/C sky130_fd_sc_hd__or3_4
XFILLER_109_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12206_ _12206_/A VGND VGND VPWR VPWR _12277_/B sky130_fd_sc_hd__inv_2
XFILLER_124_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13186_ _13186_/A _23378_/Q VGND VGND VPWR VPWR _13186_/X sky130_fd_sc_hd__or2_4
XANTENNA__22413__A _21017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19802_ _18329_/X VGND VGND VPWR VPWR _19802_/Y sky130_fd_sc_hd__inv_2
X_12137_ _12127_/B VGND VGND VPWR VPWR _12137_/Y sky130_fd_sc_hd__inv_2
X_17994_ _17928_/X _17994_/B _17994_/C VGND VGND VPWR VPWR _17994_/X sky130_fd_sc_hd__and3_4
XFILLER_123_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19733_ _19732_/Y _19730_/X _19642_/X _19730_/X VGND VGND VPWR VPWR _19733_/X sky130_fd_sc_hd__a2bb2o_4
X_12068_ _12068_/A VGND VGND VPWR VPWR _12095_/A sky130_fd_sc_hd__buf_2
X_16945_ _16938_/X _16940_/X _16942_/X _16944_/X VGND VGND VPWR VPWR _16952_/C sky130_fd_sc_hd__or4_4
XFILLER_111_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19785__B1 _19783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19664_ _19017_/X VGND VGND VPWR VPWR _19664_/X sky130_fd_sc_hd__buf_2
X_16876_ _19787_/A VGND VGND VPWR VPWR _16876_/X sky130_fd_sc_hd__buf_2
XFILLER_65_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24329__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18615_ _16622_/Y _18614_/X _16622_/Y _18614_/X VGND VGND VPWR VPWR _18615_/X sky130_fd_sc_hd__a2bb2o_4
X_15827_ _12305_/Y _15826_/X _11822_/X _15826_/X VGND VGND VPWR VPWR _24817_/D sky130_fd_sc_hd__a2bb2o_4
X_19595_ _21963_/D VGND VGND VPWR VPWR _21953_/A sky130_fd_sc_hd__inv_2
XFILLER_18_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21690__C _21646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17242__A _17242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15758_ HWDATA[8] VGND VGND VPWR VPWR _15758_/X sky130_fd_sc_hd__buf_2
X_18546_ _18541_/A _18542_/B _18546_/C VGND VGND VPWR VPWR _18546_/X sky130_fd_sc_hd__and3_4
XANTENNA__21344__B1 SSn_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14709_ _21781_/A _14703_/X _14708_/X VGND VGND VPWR VPWR _14709_/Y sky130_fd_sc_hd__a21oi_4
X_15689_ _15689_/A VGND VGND VPWR VPWR _15689_/Y sky130_fd_sc_hd__inv_2
X_18477_ _18467_/Y _18468_/Y _18477_/C VGND VGND VPWR VPWR _18478_/B sky130_fd_sc_hd__or3_4
XFILLER_127_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17428_ _17427_/Y _17425_/X _16782_/X _17425_/X VGND VGND VPWR VPWR _24317_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16771__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23964__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17359_ _17361_/B VGND VGND VPWR VPWR _17359_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20370_ _23391_/Q VGND VGND VPWR VPWR _21800_/B sky130_fd_sc_hd__inv_2
XFILLER_105_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19029_ _19029_/A VGND VGND VPWR VPWR _19029_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22040_ _22039_/X VGND VGND VPWR VPWR _22040_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23991_ _24955_/CLK _20670_/X HRESETn VGND VGND VPWR VPWR _23991_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24752__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12312__B2 _24807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22942_ _22270_/X _22939_/X _22941_/X VGND VGND VPWR VPWR _22942_/X sky130_fd_sc_hd__and3_4
XFILLER_28_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22873_ _15592_/Y _22873_/B VGND VGND VPWR VPWR _22873_/X sky130_fd_sc_hd__and2_4
X_24612_ _24612_/CLK _24612_/D HRESETn VGND VGND VPWR VPWR _24612_/Q sky130_fd_sc_hd__dfrtp_4
X_21824_ _13656_/A VGND VGND VPWR VPWR _21824_/Y sky130_fd_sc_hd__inv_2
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11823__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24543_ _24541_/CLK _24543_/D HRESETn VGND VGND VPWR VPWR _24543_/Q sky130_fd_sc_hd__dfrtp_4
X_21755_ _14752_/A _21755_/B VGND VGND VPWR VPWR _21757_/B sky130_fd_sc_hd__or2_4
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12296__A _12296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20706_ _20678_/X VGND VGND VPWR VPWR _20706_/X sky130_fd_sc_hd__buf_2
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24474_ _24649_/CLK _24474_/D HRESETn VGND VGND VPWR VPWR _16699_/A sky130_fd_sc_hd__dfrtp_4
X_21686_ _21686_/A _21816_/B VGND VGND VPWR VPWR _21686_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__16762__B1 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12379__B2 _24810_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23425_ _23682_/CLK _23425_/D VGND VGND VPWR VPWR _23425_/Q sky130_fd_sc_hd__dfxtp_4
X_20637_ _20637_/A VGND VGND VPWR VPWR _20637_/Y sky130_fd_sc_hd__inv_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25540__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16514__B1 _16340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23356_ _23343_/X VGND VGND VPWR VPWR IRQ[2] sky130_fd_sc_hd__buf_2
X_20568_ _14428_/Y _20556_/X _20547_/X _20567_/X VGND VGND VPWR VPWR _20569_/A sky130_fd_sc_hd__a211o_4
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22307_ _22306_/Y _21336_/A _14405_/Y _21338_/X VGND VGND VPWR VPWR _22308_/A sky130_fd_sc_hd__o22a_4
X_23287_ _23119_/X _23285_/X _23121_/X _23286_/X VGND VGND VPWR VPWR _23288_/B sky130_fd_sc_hd__o22a_4
X_20499_ _23996_/Q _20512_/B _20459_/X VGND VGND VPWR VPWR _20499_/X sky130_fd_sc_hd__a21o_4
XANTENNA__14242__A1_N _14241_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13040_ _13026_/A _13037_/B _13039_/X VGND VGND VPWR VPWR _13041_/A sky130_fd_sc_hd__or3_4
X_25026_ _25020_/CLK _15170_/X HRESETn VGND VGND VPWR VPWR _25026_/Q sky130_fd_sc_hd__dfrtp_4
X_22238_ _22246_/A _22238_/B VGND VGND VPWR VPWR _22238_/X sky130_fd_sc_hd__or2_4
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22169_ _12109_/Y _12097_/X _18374_/Y _12071_/A VGND VGND VPWR VPWR _22169_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16231__A _11803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14991_ _14991_/A VGND VGND VPWR VPWR _14991_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24493__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13500__B1 _11829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19767__B1 _19721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13942_ _13919_/X _13920_/X _13942_/C _13958_/C VGND VGND VPWR VPWR _13951_/A sky130_fd_sc_hd__or4_4
X_16730_ _16730_/A VGND VGND VPWR VPWR _16730_/X sky130_fd_sc_hd__buf_2
XFILLER_8_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24422__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12597__A2_N _12514_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16661_ _16660_/Y _16658_/X _16393_/X _16658_/X VGND VGND VPWR VPWR _16661_/X sky130_fd_sc_hd__a2bb2o_4
X_13873_ _13871_/X _13872_/X _14263_/A _13867_/X VGND VGND VPWR VPWR _25236_/D sky130_fd_sc_hd__o22a_4
XFILLER_62_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22118__A2 _22101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15612_ _15561_/X VGND VGND VPWR VPWR _15612_/X sky130_fd_sc_hd__buf_2
X_18400_ _18400_/A VGND VGND VPWR VPWR _18400_/Y sky130_fd_sc_hd__inv_2
X_12824_ _24794_/Q VGND VGND VPWR VPWR _12824_/Y sky130_fd_sc_hd__inv_2
X_16592_ _16592_/A VGND VGND VPWR VPWR _16592_/Y sky130_fd_sc_hd__inv_2
X_19380_ _19376_/Y _19379_/X _19313_/X _19379_/X VGND VGND VPWR VPWR _23748_/D sky130_fd_sc_hd__a2bb2o_4
X_15543_ _15542_/Y _15538_/X HADDR[0] _15538_/X VGND VGND VPWR VPWR _24912_/D sky130_fd_sc_hd__a2bb2o_4
X_18331_ _24196_/Q VGND VGND VPWR VPWR _18331_/X sky130_fd_sc_hd__buf_2
X_12755_ _22546_/A VGND VGND VPWR VPWR _12755_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11814__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11706_/A VGND VGND VPWR VPWR _11706_/Y sky130_fd_sc_hd__inv_2
X_18262_ _18262_/A VGND VGND VPWR VPWR _18262_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _16359_/A VGND VGND VPWR VPWR _15474_/X sky130_fd_sc_hd__buf_2
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12686_/A _12686_/B _12685_/Y VGND VGND VPWR VPWR _25404_/D sky130_fd_sc_hd__and3_4
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _25127_/Q VGND VGND VPWR VPWR _14425_/Y sky130_fd_sc_hd__inv_2
X_17213_ _16305_/Y _17237_/A _16305_/Y _17237_/A VGND VGND VPWR VPWR _17213_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21312__A _21019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18193_ _18097_/A _18185_/X _18192_/X VGND VGND VPWR VPWR _18193_/X sky130_fd_sc_hd__and3_4
XFILLER_50_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25281__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22127__B _22124_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_106_0_HCLK clkbuf_7_53_0_HCLK/X VGND VGND VPWR VPWR _24330_/CLK sky130_fd_sc_hd__clkbuf_1
X_17144_ _17038_/C _17148_/A VGND VGND VPWR VPWR _17145_/C sky130_fd_sc_hd__nand2_4
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _14344_/X VGND VGND VPWR VPWR _14356_/X sky130_fd_sc_hd__buf_2
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16505__B1 _16231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_169_0_HCLK clkbuf_7_84_0_HCLK/X VGND VGND VPWR VPWR _23714_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22841__A3 _16728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13307_ _13269_/A _23375_/Q VGND VGND VPWR VPWR _13309_/B sky130_fd_sc_hd__or2_4
X_17075_ _17384_/B _17071_/B _17075_/C VGND VGND VPWR VPWR _17076_/A sky130_fd_sc_hd__or3_4
X_14287_ _13522_/A VGND VGND VPWR VPWR _14291_/A sky130_fd_sc_hd__inv_2
X_16026_ _24722_/Q VGND VGND VPWR VPWR _16026_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13238_ _13386_/A _13238_/B _13238_/C VGND VGND VPWR VPWR _13244_/B sky130_fd_sc_hd__and3_4
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13169_ _13251_/A VGND VGND VPWR VPWR _18344_/A sky130_fd_sc_hd__buf_2
XFILLER_97_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18273__A3 _11867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17977_ _18104_/A _23451_/Q VGND VGND VPWR VPWR _17978_/C sky130_fd_sc_hd__or2_4
XANTENNA__15492__B1 HWRITE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19716_ _19714_/Y _19712_/X _19715_/X _19712_/X VGND VGND VPWR VPWR _23633_/D sky130_fd_sc_hd__a2bb2o_4
X_16928_ _24250_/Q VGND VGND VPWR VPWR _16928_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19647_ _19644_/Y _19639_/X _19645_/X _19646_/X VGND VGND VPWR VPWR _23658_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18430__B1 _16230_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16859_ _16880_/A VGND VGND VPWR VPWR _16859_/X sky130_fd_sc_hd__buf_2
XANTENNA__15244__B1 _15199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19578_ _23677_/Q VGND VGND VPWR VPWR _21176_/B sky130_fd_sc_hd__inv_2
XFILLER_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18529_ _18524_/A _18523_/X _18498_/X _18525_/Y VGND VGND VPWR VPWR _18530_/A sky130_fd_sc_hd__a211o_4
XANTENNA__21868__A1 _16156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21868__B2 _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25369__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13005__A _12294_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21540_ _14487_/Y _14258_/A VGND VGND VPWR VPWR _21540_/X sky130_fd_sc_hd__or2_4
XANTENNA__16744__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11744__A2_N _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22817__B1 _21050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16961__A1_N _24709_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21471_ _18293_/B VGND VGND VPWR VPWR _21477_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_65_0_HCLK clkbuf_6_32_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_65_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16316__A _16288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23210_ _23210_/A _23269_/B VGND VGND VPWR VPWR _23210_/X sky130_fd_sc_hd__or2_4
X_20422_ _14380_/B VGND VGND VPWR VPWR _20422_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12230__B1 _12278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24190_ _23377_/CLK _24190_/D HRESETn VGND VGND VPWR VPWR _24190_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23141_ _22466_/A VGND VGND VPWR VPWR _23141_/X sky130_fd_sc_hd__buf_2
X_20353_ _21654_/B _20352_/X _19629_/A _20352_/X VGND VGND VPWR VPWR _20353_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23965__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12282__C _12282_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20284_ _22006_/B _20278_/X _19981_/X _20283_/X VGND VGND VPWR VPWR _23425_/D sky130_fd_sc_hd__a2bb2o_4
X_23072_ _23072_/A _21017_/B VGND VGND VPWR VPWR _23075_/B sky130_fd_sc_hd__or2_4
XANTENNA__24933__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22023_ _21664_/A _22023_/B VGND VGND VPWR VPWR _22023_/X sky130_fd_sc_hd__or2_4
XFILLER_103_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16051__A _24712_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_25_0_HCLK_A clkbuf_4_12_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23974_ _24943_/CLK _20632_/Y HRESETn VGND VGND VPWR VPWR _20629_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_112_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22925_ _24521_/Q _22922_/X _22923_/X _22924_/X VGND VGND VPWR VPWR _22926_/C sky130_fd_sc_hd__a211o_4
XFILLER_17_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22856_ _22763_/A _22856_/B VGND VGND VPWR VPWR _22856_/X sky130_fd_sc_hd__and2_4
XFILLER_45_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21807_ _21477_/A _21807_/B VGND VGND VPWR VPWR _21807_/X sky130_fd_sc_hd__or2_4
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22787_ _22787_/A _22873_/B VGND VGND VPWR VPWR _22787_/X sky130_fd_sc_hd__and2_4
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19921__B1 _19790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12540_ _25412_/Q _12539_/A _12656_/A _12539_/Y VGND VGND VPWR VPWR _12540_/X sky130_fd_sc_hd__o22a_4
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24526_ _24557_/CLK _16564_/X HRESETn VGND VGND VPWR VPWR _24526_/Q sky130_fd_sc_hd__dfrtp_4
X_21738_ _16711_/Y _21582_/B VGND VGND VPWR VPWR _21738_/X sky130_fd_sc_hd__and2_4
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16735__B1 _16380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25039__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12471_ _12209_/Y _12269_/Y _12278_/B _12471_/D VGND VGND VPWR VPWR _12471_/X sky130_fd_sc_hd__or4_4
X_24457_ _24457_/CLK _24457_/D HRESETn VGND VGND VPWR VPWR _24457_/Q sky130_fd_sc_hd__dfrtp_4
X_21669_ _21477_/A _21669_/B VGND VGND VPWR VPWR _21671_/B sky130_fd_sc_hd__or2_4
X_14210_ _20657_/A _14210_/B VGND VGND VPWR VPWR _14210_/X sky130_fd_sc_hd__or2_4
XFILLER_71_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23408_ _24209_/CLK _20328_/X VGND VGND VPWR VPWR _23408_/Q sky130_fd_sc_hd__dfxtp_4
X_15190_ _15190_/A _15185_/Y _15189_/X VGND VGND VPWR VPWR _15191_/A sky130_fd_sc_hd__or3_4
X_24388_ _24362_/CLK _24388_/D HRESETn VGND VGND VPWR VPWR _24388_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14141_ _23949_/D _14140_/Y _25128_/Q _23949_/D VGND VGND VPWR VPWR _25208_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19537__A _16725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23339_ _18265_/Y _24198_/Q _17480_/Y _24209_/Q VGND VGND VPWR VPWR _23339_/X sky130_fd_sc_hd__a2bb2o_4
X_14072_ _14036_/C _14071_/X VGND VGND VPWR VPWR _14073_/B sky130_fd_sc_hd__nor2_4
XANTENNA__15784__B _15784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13023_ _13023_/A _13023_/B VGND VGND VPWR VPWR _13024_/C sky130_fd_sc_hd__or2_4
X_17900_ _17900_/A _17900_/B VGND VGND VPWR VPWR _17900_/X sky130_fd_sc_hd__and2_4
XANTENNA__24674__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25009_ _25010_/CLK _25009_/D HRESETn VGND VGND VPWR VPWR _25009_/Q sky130_fd_sc_hd__dfrtp_4
X_18880_ _23942_/Q _18879_/X VGND VGND VPWR VPWR _18880_/X sky130_fd_sc_hd__or2_4
XFILLER_126_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22898__A _21525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24603__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17831_ _17833_/B VGND VGND VPWR VPWR _17831_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17762_ _17762_/A _17761_/X VGND VGND VPWR VPWR _17762_/X sky130_fd_sc_hd__or2_4
X_14974_ _14965_/X _14974_/B _14970_/X _14973_/X VGND VGND VPWR VPWR _14984_/C sky130_fd_sc_hd__or4_4
XFILLER_43_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22410__B _21073_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19501_ _22004_/B _19495_/X _11939_/X _19500_/X VGND VGND VPWR VPWR _23706_/D sky130_fd_sc_hd__a2bb2o_4
X_16713_ _16711_/Y _16707_/X _16359_/X _16712_/X VGND VGND VPWR VPWR _16713_/X sky130_fd_sc_hd__a2bb2o_4
X_13925_ _24958_/Q VGND VGND VPWR VPWR _13956_/A sky130_fd_sc_hd__buf_2
X_17693_ _17662_/B _17688_/X VGND VGND VPWR VPWR _17694_/B sky130_fd_sc_hd__nand2_4
XANTENNA__20211__A _20210_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23225__C _22132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19432_ _19430_/Y _19425_/X _19407_/X _19431_/X VGND VGND VPWR VPWR _19432_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11833__A _13835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13856_ _23989_/Q VGND VGND VPWR VPWR _13856_/Y sky130_fd_sc_hd__inv_2
X_16644_ _16643_/Y VGND VGND VPWR VPWR _16645_/A sky130_fd_sc_hd__buf_2
XFILLER_78_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21026__B _21026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12807_ _22660_/A _22651_/A _22660_/A _22651_/A VGND VGND VPWR VPWR _12807_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19363_ _23753_/Q VGND VGND VPWR VPWR _19363_/Y sky130_fd_sc_hd__inv_2
X_13787_ _13787_/A VGND VGND VPWR VPWR _15662_/A sky130_fd_sc_hd__buf_2
X_16575_ _16558_/A VGND VGND VPWR VPWR _16575_/X sky130_fd_sc_hd__buf_2
XFILLER_16_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13470__D _12059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25462__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19912__B1 _19777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18314_ _18314_/A VGND VGND VPWR VPWR _18314_/Y sky130_fd_sc_hd__inv_2
X_12738_ _12529_/Y _12629_/X _12648_/A _12736_/B VGND VGND VPWR VPWR _12739_/A sky130_fd_sc_hd__a211o_4
X_15526_ _24920_/Q VGND VGND VPWR VPWR _15526_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19294_ _18996_/X VGND VGND VPWR VPWR _19294_/X sky130_fd_sc_hd__buf_2
XANTENNA__16726__B1 _16720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15457_ _13897_/X _20602_/A _15446_/A _13895_/X _15452_/X VGND VGND VPWR VPWR _15457_/X
+ sky130_fd_sc_hd__a32o_4
X_18245_ _18235_/X _18237_/X _16600_/X _22507_/A _18238_/X VGND VGND VPWR VPWR _24222_/D
+ sky130_fd_sc_hd__a32o_4
X_12669_ _25409_/Q _12669_/B VGND VGND VPWR VPWR _12669_/X sky130_fd_sc_hd__or2_4
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14408_ _11733_/A _14475_/B VGND VGND VPWR VPWR _14408_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15040__A _15034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15388_ _15159_/X _15388_/B _15388_/C _15421_/A VGND VGND VPWR VPWR _15388_/X sky130_fd_sc_hd__or4_4
X_18176_ _18176_/A _18174_/X _18176_/C VGND VGND VPWR VPWR _18177_/C sky130_fd_sc_hd__and3_4
XFILLER_102_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14339_ _14339_/A VGND VGND VPWR VPWR _14339_/Y sky130_fd_sc_hd__inv_2
X_17127_ _17023_/Y _17043_/Y VGND VGND VPWR VPWR _17161_/A sky130_fd_sc_hd__or2_4
XFILLER_7_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17058_ _17057_/X VGND VGND VPWR VPWR _17058_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23224__B1 _25383_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16009_ _24729_/Q VGND VGND VPWR VPWR _16009_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13495__A _16183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_HCLK clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__24344__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18651__B1 _16585_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21862__D _21861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20971_ _14181_/B _20970_/X _20978_/B VGND VGND VPWR VPWR _23950_/D sky130_fd_sc_hd__o21a_4
XFILLER_122_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15217__B1 _15199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17014__A1_N _24731_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11743__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22710_ _23306_/A _22706_/X _22710_/C VGND VGND VPWR VPWR _22710_/X sky130_fd_sc_hd__and3_4
X_23690_ _23384_/CLK _19545_/X VGND VGND VPWR VPWR _23690_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22641_ _22625_/Y _22630_/Y _22638_/Y _21437_/X _22640_/X VGND VGND VPWR VPWR _22642_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_22_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25360_ _25330_/CLK _12967_/X HRESETn VGND VGND VPWR VPWR _25360_/Q sky130_fd_sc_hd__dfrtp_4
X_22572_ _24444_/Q _22525_/X _22526_/X VGND VGND VPWR VPWR _22572_/X sky130_fd_sc_hd__o21a_4
X_24311_ _24187_/CLK _24311_/D HRESETn VGND VGND VPWR VPWR _24311_/Q sky130_fd_sc_hd__dfstp_4
X_21523_ _15784_/B VGND VGND VPWR VPWR _22489_/A sky130_fd_sc_hd__buf_2
X_25291_ _25290_/CLK _25291_/D HRESETn VGND VGND VPWR VPWR _13532_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16046__A _24714_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24242_ _24186_/CLK _17908_/X HRESETn VGND VGND VPWR VPWR _17893_/A sky130_fd_sc_hd__dfrtp_4
X_21454_ _21454_/A VGND VGND VPWR VPWR _21460_/A sky130_fd_sc_hd__buf_2
X_20405_ _20399_/Y VGND VGND VPWR VPWR _20405_/X sky130_fd_sc_hd__buf_2
XFILLER_119_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24173_ _25029_/CLK _24173_/D HRESETn VGND VGND VPWR VPWR _18438_/A sky130_fd_sc_hd__dfrtp_4
X_21385_ _21385_/A _21385_/B VGND VGND VPWR VPWR _21386_/C sky130_fd_sc_hd__or2_4
XANTENNA__18261__A _18261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_152_0_HCLK clkbuf_7_76_0_HCLK/X VGND VGND VPWR VPWR _24187_/CLK sky130_fd_sc_hd__clkbuf_1
X_23124_ _23124_/A _23124_/B VGND VGND VPWR VPWR _23124_/Y sky130_fd_sc_hd__nor2_4
X_20336_ _20335_/Y _20326_/Y _19771_/X _20326_/Y VGND VGND VPWR VPWR _23404_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23055_ _20779_/Y _22988_/X _20918_/Y _21211_/X VGND VGND VPWR VPWR _23055_/X sky130_fd_sc_hd__o22a_4
X_20267_ _21626_/B _20266_/X _16879_/A _20266_/X VGND VGND VPWR VPWR _20267_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21777__B1 _21821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24085__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22006_ _22005_/X _22006_/B VGND VGND VPWR VPWR _22006_/X sky130_fd_sc_hd__or2_4
XANTENNA__18642__B1 _16611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20198_ _20198_/A VGND VGND VPWR VPWR _21882_/B sky130_fd_sc_hd__inv_2
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24014__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11971_ _11969_/Y _11970_/X _11967_/X VGND VGND VPWR VPWR _11971_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_29_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23957_ _24070_/CLK _25171_/Q HRESETn VGND VGND VPWR VPWR _23957_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12749__A _12749_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13710_ _13690_/A _13689_/X VGND VGND VPWR VPWR _13710_/Y sky130_fd_sc_hd__nand2_4
XFILLER_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22908_ _22419_/X VGND VGND VPWR VPWR _22908_/X sky130_fd_sc_hd__buf_2
X_14690_ _13748_/A _14752_/A _13748_/A _14752_/A VGND VGND VPWR VPWR _14719_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23888_ _23887_/CLK _18979_/X VGND VGND VPWR VPWR _18976_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12468__B _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20752__B2 _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13641_ _12026_/X _13524_/B _13527_/B VGND VGND VPWR VPWR _13642_/B sky130_fd_sc_hd__o21a_4
XANTENNA__23342__A _23342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22839_ _22819_/X _22823_/Y _22830_/Y _22838_/X VGND VGND VPWR VPWR _22852_/C sky130_fd_sc_hd__a211o_4
XFILLER_38_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14431__B2 _14408_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16360_ _16358_/Y _16356_/X _16359_/X _16356_/X VGND VGND VPWR VPWR _24602_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17340__A _22659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _25245_/Q VGND VGND VPWR VPWR _13572_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16708__B1 _16528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15779__B _15674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15311_ _15313_/B VGND VGND VPWR VPWR _15312_/B sky130_fd_sc_hd__inv_2
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _24852_/Q VGND VGND VPWR VPWR _12523_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24509_ _24553_/CLK _16607_/X HRESETn VGND VGND VPWR VPWR _24509_/Q sky130_fd_sc_hd__dfrtp_4
X_16291_ _24627_/Q VGND VGND VPWR VPWR _16291_/Y sky130_fd_sc_hd__inv_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25489_ _25488_/CLK _25489_/D HRESETn VGND VGND VPWR VPWR _11702_/C sky130_fd_sc_hd__dfrtp_4
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15242_ _15209_/A _15240_/A VGND VGND VPWR VPWR _15242_/X sky130_fd_sc_hd__or2_4
X_18030_ _18104_/A _20216_/A VGND VGND VPWR VPWR _18031_/C sky130_fd_sc_hd__or2_4
X_12454_ _12248_/A _12454_/B VGND VGND VPWR VPWR _12454_/X sky130_fd_sc_hd__or2_4
XANTENNA__24855__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15173_ _15180_/A _15166_/B _15172_/X VGND VGND VPWR VPWR _15173_/X sky130_fd_sc_hd__or3_4
XANTENNA__15795__A _15795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12385_ _12385_/A _12385_/B _12266_/Y _12397_/B VGND VGND VPWR VPWR _12385_/X sky130_fd_sc_hd__or4_4
XANTENNA__18171__A _18024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14124_ _14124_/A VGND VGND VPWR VPWR _14125_/A sky130_fd_sc_hd__buf_2
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23206__B1 _22997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19981_ _11932_/A VGND VGND VPWR VPWR _19981_/X sky130_fd_sc_hd__buf_2
XFILLER_125_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14055_ _20531_/A _13976_/X _14052_/X _14054_/Y VGND VGND VPWR VPWR _14056_/A sky130_fd_sc_hd__o22a_4
X_18932_ _13310_/B VGND VGND VPWR VPWR _18932_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13006_ _13038_/A _13004_/X _13005_/X VGND VGND VPWR VPWR _13006_/X sky130_fd_sc_hd__and3_4
XFILLER_84_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18863_ _24560_/Q _18672_/Y _24554_/Q _18656_/Y VGND VGND VPWR VPWR _18864_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22421__A _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21705__A2_N _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17814_ _16900_/Y _17814_/B VGND VGND VPWR VPWR _17815_/C sky130_fd_sc_hd__or2_4
X_18794_ _18794_/A VGND VGND VPWR VPWR _18794_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17745_ _17745_/A VGND VGND VPWR VPWR _17747_/C sky130_fd_sc_hd__inv_2
X_14957_ _15193_/A _24424_/Q _14955_/Y _24424_/Q VGND VGND VPWR VPWR _14963_/B sky130_fd_sc_hd__a2bb2o_4
X_13908_ _13905_/X _13908_/B VGND VGND VPWR VPWR _13908_/X sky130_fd_sc_hd__or2_4
XFILLER_130_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19730__A _19729_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17676_ _17676_/A _17676_/B VGND VGND VPWR VPWR _17677_/C sky130_fd_sc_hd__nand2_4
X_14888_ _25026_/Q VGND VGND VPWR VPWR _14888_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21940__B1 _17722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19415_ _19401_/A VGND VGND VPWR VPWR _19415_/X sky130_fd_sc_hd__buf_2
X_16627_ _13743_/B _16172_/B _16634_/B VGND VGND VPWR VPWR _16627_/X sky130_fd_sc_hd__a21o_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13839_ _13821_/A VGND VGND VPWR VPWR _13839_/X sky130_fd_sc_hd__buf_2
XFILLER_56_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19346_ _19333_/Y VGND VGND VPWR VPWR _19346_/X sky130_fd_sc_hd__buf_2
XANTENNA__22496__A1 _16599_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16558_ _16558_/A VGND VGND VPWR VPWR _16558_/X sky130_fd_sc_hd__buf_2
XFILLER_52_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15509_ _15508_/Y _15504_/X HADDR[15] _15504_/X VGND VGND VPWR VPWR _15509_/X sky130_fd_sc_hd__a2bb2o_4
X_19277_ _23783_/Q VGND VGND VPWR VPWR _21607_/B sky130_fd_sc_hd__inv_2
X_16489_ _16488_/Y _16486_/X _16403_/X _16486_/X VGND VGND VPWR VPWR _24554_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18228_ _13815_/X VGND VGND VPWR VPWR _18230_/A sky130_fd_sc_hd__buf_2
XANTENNA__22799__A2 _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24596__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18159_ _18191_/A _18159_/B _18158_/X VGND VGND VPWR VPWR _18159_/X sky130_fd_sc_hd__and3_4
XFILLER_89_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24525__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21170_ _21186_/A _21170_/B _21169_/X VGND VGND VPWR VPWR _21170_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_225_0_HCLK clkbuf_8_225_0_HCLK/A VGND VGND VPWR VPWR _24785_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12841__B _12841_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20121_ _21385_/B _20118_/X _20099_/X _20118_/X VGND VGND VPWR VPWR _20121_/X sky130_fd_sc_hd__a2bb2o_4
X_20052_ _23513_/Q VGND VGND VPWR VPWR _21904_/B sky130_fd_sc_hd__inv_2
XFILLER_98_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24860_ _24847_/CLK _24860_/D HRESETn VGND VGND VPWR VPWR _12555_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23146__B _23145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23811_ _23818_/CLK _23811_/D VGND VGND VPWR VPWR _19200_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_22_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24791_ _24800_/CLK _15883_/X HRESETn VGND VGND VPWR VPWR _22895_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25384__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22723__A2 _22525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23742_ _23446_/CLK _23742_/D VGND VGND VPWR VPWR _18165_/B sky130_fd_sc_hd__dfxtp_4
X_20954_ _12001_/A _20955_/B VGND VGND VPWR VPWR _20954_/X sky130_fd_sc_hd__and2_4
XFILLER_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16938__B1 _22556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25313__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _23689_/CLK _19596_/X VGND VGND VPWR VPWR _21963_/D sky130_fd_sc_hd__dfxtp_4
X_20885_ _24044_/Q _20879_/X _20884_/Y VGND VGND VPWR VPWR _20885_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15610__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23279__A3 _22127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25412_ _25400_/CLK _12657_/X HRESETn VGND VGND VPWR VPWR _25412_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22624_ _21040_/A _22623_/X _22396_/C _24854_/Q _22547_/X VGND VGND VPWR VPWR _22625_/B
+ sky130_fd_sc_hd__a32o_4
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25343_ _23370_/CLK _13049_/X HRESETn VGND VGND VPWR VPWR _25343_/Q sky130_fd_sc_hd__dfrtp_4
X_22555_ _21064_/A _22552_/X _21098_/X _22554_/X VGND VGND VPWR VPWR _22555_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__17363__B1 _17289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21506_ _21505_/X VGND VGND VPWR VPWR _21506_/Y sky130_fd_sc_hd__inv_2
X_25274_ _24252_/CLK _25274_/D HRESETn VGND VGND VPWR VPWR _25274_/Q sky130_fd_sc_hd__dfrtp_4
X_22486_ _15791_/A _22484_/X _22485_/X _11824_/A _22915_/A VGND VGND VPWR VPWR _22486_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12304__A2_N _24823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_35_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_71_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24225_ _24715_/CLK _18241_/X HRESETn VGND VGND VPWR VPWR _24225_/Q sky130_fd_sc_hd__dfrtp_4
X_21437_ _21024_/X VGND VGND VPWR VPWR _21437_/X sky130_fd_sc_hd__buf_2
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24266__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12170_ _12159_/X _12169_/X SCLK_S3 _12159_/X VGND VGND VPWR VPWR _12170_/X sky130_fd_sc_hd__a2bb2o_4
X_24156_ _24151_/CLK _18568_/X HRESETn VGND VGND VPWR VPWR _24156_/Q sky130_fd_sc_hd__dfrtp_4
X_21368_ _21368_/A _22575_/A VGND VGND VPWR VPWR _21368_/X sky130_fd_sc_hd__and2_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18863__B1 _24554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23107_ _24624_/Q _22898_/X VGND VGND VPWR VPWR _23107_/X sky130_fd_sc_hd__or2_4
X_20319_ _20318_/X VGND VGND VPWR VPWR _22389_/B sky130_fd_sc_hd__buf_2
X_24087_ _25301_/CLK _24087_/D HRESETn VGND VGND VPWR VPWR _24087_/Q sky130_fd_sc_hd__dfrtp_4
X_21299_ _23097_/A VGND VGND VPWR VPWR _21299_/X sky130_fd_sc_hd__buf_2
XANTENNA__17038__C _17038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17536__A1_N _11798_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18615__B1 _16622_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22411__A1 _21413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23038_ _22897_/A _23037_/X VGND VGND VPWR VPWR _23038_/X sky130_fd_sc_hd__and2_4
XFILLER_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22241__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15860_ _23035_/A VGND VGND VPWR VPWR _21026_/B sky130_fd_sc_hd__buf_2
XFILLER_114_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14811_ _14809_/A VGND VGND VPWR VPWR _14811_/X sky130_fd_sc_hd__buf_2
X_15791_ _15791_/A _15925_/B VGND VGND VPWR VPWR _15817_/A sky130_fd_sc_hd__or2_4
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24989_ _24984_/CLK _24989_/D HRESETn VGND VGND VPWR VPWR _24989_/Q sky130_fd_sc_hd__dfrtp_4
X_17530_ _11811_/Y _17571_/A _11811_/Y _17571_/A VGND VGND VPWR VPWR _17530_/X sky130_fd_sc_hd__a2bb2o_4
X_11954_ _19885_/A VGND VGND VPWR VPWR _11954_/Y sky130_fd_sc_hd__inv_2
X_14742_ _22038_/A VGND VGND VPWR VPWR _14742_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21922__B1 _17722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25054__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23072__A _23072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14673_ _13613_/X _13633_/B _14671_/X VGND VGND VPWR VPWR _14673_/X sky130_fd_sc_hd__o21a_4
X_17461_ _17458_/X _17489_/A VGND VGND VPWR VPWR _17461_/X sky130_fd_sc_hd__or2_4
X_11885_ _13678_/B _11884_/X _11870_/A _11872_/X VGND VGND VPWR VPWR _11886_/A sky130_fd_sc_hd__a211o_4
XFILLER_60_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19200_ _19200_/A VGND VGND VPWR VPWR _19200_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15601__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13624_ _13624_/A VGND VGND VPWR VPWR _14658_/A sky130_fd_sc_hd__inv_2
X_16412_ _24583_/Q VGND VGND VPWR VPWR _16412_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_117_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_235_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17392_ _20629_/A _20625_/A VGND VGND VPWR VPWR _17392_/X sky130_fd_sc_hd__or2_4
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19131_ _19126_/Y _19130_/X _19018_/X _19130_/X VGND VGND VPWR VPWR _23836_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20489__B1 _20481_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13555_ _25257_/Q VGND VGND VPWR VPWR _22726_/A sky130_fd_sc_hd__inv_2
X_16343_ _16324_/A VGND VGND VPWR VPWR _16343_/X sky130_fd_sc_hd__buf_2
XFILLER_41_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12506_ _13008_/B VGND VGND VPWR VPWR _13042_/A sky130_fd_sc_hd__buf_2
X_16274_ _15655_/X _15993_/Y _16270_/X _24632_/Q _16273_/X VGND VGND VPWR VPWR _16274_/X
+ sky130_fd_sc_hd__a32o_4
X_19062_ _19062_/A VGND VGND VPWR VPWR _19062_/Y sky130_fd_sc_hd__inv_2
X_13486_ _25307_/Q VGND VGND VPWR VPWR _13486_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15225_ _15216_/A _15219_/X _15225_/C VGND VGND VPWR VPWR _15225_/X sky130_fd_sc_hd__and3_4
X_18013_ _17929_/A _19178_/A VGND VGND VPWR VPWR _18013_/X sky130_fd_sc_hd__or2_4
XFILLER_16_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21320__A _23170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12437_ _12429_/X _12435_/X _12436_/X VGND VGND VPWR VPWR _25441_/D sky130_fd_sc_hd__and3_4
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12942__A _12819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15156_ _15155_/Y _16378_/A _15155_/Y _16378_/A VGND VGND VPWR VPWR _15161_/B sky130_fd_sc_hd__a2bb2o_4
X_12368_ _12368_/A VGND VGND VPWR VPWR _12368_/Y sky130_fd_sc_hd__inv_2
X_14107_ _14381_/A _14096_/X _14107_/C VGND VGND VPWR VPWR _14108_/A sky130_fd_sc_hd__or3_4
XANTENNA__20661__B1 _17387_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15087_ _24989_/Q VGND VGND VPWR VPWR _15087_/Y sky130_fd_sc_hd__inv_2
X_19964_ _19964_/A VGND VGND VPWR VPWR _19964_/X sky130_fd_sc_hd__buf_2
XFILLER_99_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12299_ _12299_/A VGND VGND VPWR VPWR _12299_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14038_ _14037_/X VGND VGND VPWR VPWR _14038_/Y sky130_fd_sc_hd__inv_2
X_18915_ _18913_/Y _18914_/X _16885_/X _18914_/X VGND VGND VPWR VPWR _23911_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18606__B1 _16581_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23989__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19895_ _19902_/A VGND VGND VPWR VPWR _19895_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_55_0_HCLK clkbuf_8_55_0_HCLK/A VGND VGND VPWR VPWR _24391_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20413__B1 _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17245__A _17244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18846_ _16495_/Y _24130_/Q _16485_/A _18749_/A VGND VGND VPWR VPWR _18849_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23918__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18777_ _18759_/A _18775_/X _18776_/X VGND VGND VPWR VPWR _18777_/X sky130_fd_sc_hd__and3_4
X_15989_ _15788_/X _15857_/A _15927_/X _24735_/Q _15933_/A VGND VGND VPWR VPWR _24735_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22166__B1 _25426_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17728_ _17728_/A VGND VGND VPWR VPWR _21491_/A sky130_fd_sc_hd__buf_2
XANTENNA__19031__B1 _18961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17659_ _17571_/Y _17653_/X _17656_/B _17590_/X VGND VGND VPWR VPWR _17660_/A sky130_fd_sc_hd__a211o_4
XFILLER_91_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20670_ _20665_/X _20669_/X _20602_/X VGND VGND VPWR VPWR _20670_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21214__B _21859_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24777__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19329_ _23765_/Q VGND VGND VPWR VPWR _19329_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21141__B2 _14433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24706__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22340_ _22005_/X _22340_/B VGND VGND VPWR VPWR _22340_/X sky130_fd_sc_hd__or2_4
XFILLER_137_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22326__A _21458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22271_ _21700_/X VGND VGND VPWR VPWR _22271_/X sky130_fd_sc_hd__buf_2
XFILLER_117_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14770__C _14555_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24010_ _24041_/CLK _20737_/X HRESETn VGND VGND VPWR VPWR _13133_/A sky130_fd_sc_hd__dfrtp_4
X_21222_ _14679_/A VGND VGND VPWR VPWR _21252_/A sky130_fd_sc_hd__buf_2
XFILLER_89_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18845__B1 _24544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21153_ _16268_/Y _21556_/A _16449_/A _21152_/X VGND VGND VPWR VPWR _21159_/B sky130_fd_sc_hd__a211o_4
XFILLER_137_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20104_ _19844_/X _13748_/X VGND VGND VPWR VPWR _20105_/A sky130_fd_sc_hd__and2_4
XANTENNA__22699__C _21859_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21084_ _21071_/A VGND VGND VPWR VPWR _21085_/A sky130_fd_sc_hd__buf_2
XFILLER_8_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20035_ _20035_/A VGND VGND VPWR VPWR _20035_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24912_ _24923_/CLK _24912_/D HRESETn VGND VGND VPWR VPWR _15542_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12893__B1 _12874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24843_ _24847_/CLK _24843_/D HRESETn VGND VGND VPWR VPWR _12562_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_67_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15831__B1 _15620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19370__A _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24774_ _24780_/CLK _24774_/D HRESETn VGND VGND VPWR VPWR _24774_/Q sky130_fd_sc_hd__dfrtp_4
X_21986_ _17893_/A _21985_/B VGND VGND VPWR VPWR _21987_/C sky130_fd_sc_hd__or2_4
XPHY_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _23722_/CLK _19443_/X VGND VGND VPWR VPWR _18204_/B sky130_fd_sc_hd__dfxtp_4
X_20937_ _20936_/X VGND VGND VPWR VPWR _20937_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14398__B1 _14239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11669_/Y _24216_/Q _11669_/Y _24216_/Q VGND VGND VPWR VPWR _11670_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23656_ _24197_/CLK _23656_/D VGND VGND VPWR VPWR _13356_/B sky130_fd_sc_hd__dfxtp_4
X_20868_ _20867_/Y _20861_/Y _13662_/B VGND VGND VPWR VPWR _20868_/X sky130_fd_sc_hd__o21a_4
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22607_ _22574_/X _22582_/Y _22586_/X _22607_/D VGND VGND VPWR VPWR HRDATA[11] sky130_fd_sc_hd__or4_4
XANTENNA__21722__A1_N _16261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23587_ _23516_/CLK _23587_/D VGND VGND VPWR VPWR _23587_/Q sky130_fd_sc_hd__dfxtp_4
X_20799_ _20799_/A VGND VGND VPWR VPWR _20799_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12243__A2_N _24748_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24447__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13340_ _13303_/A _13340_/B VGND VGND VPWR VPWR _13340_/X sky130_fd_sc_hd__or2_4
X_25326_ _25351_/CLK _13105_/Y HRESETn VGND VGND VPWR VPWR _25326_/Q sky130_fd_sc_hd__dfrtp_4
X_22538_ _22537_/X VGND VGND VPWR VPWR _22538_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15898__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13271_ _13309_/A _13271_/B _13270_/X VGND VGND VPWR VPWR _13271_/X sky130_fd_sc_hd__and3_4
X_25257_ _24720_/CLK _25257_/D HRESETn VGND VGND VPWR VPWR _25257_/Q sky130_fd_sc_hd__dfrtp_4
X_22469_ _22763_/A _22468_/X VGND VGND VPWR VPWR _22488_/B sky130_fd_sc_hd__and2_4
X_15010_ _24435_/Q VGND VGND VPWR VPWR _15010_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12222_ _25429_/Q _22465_/A _12220_/X _12221_/Y VGND VGND VPWR VPWR _12222_/X sky130_fd_sc_hd__o22a_4
X_24208_ _24208_/CLK _18269_/X HRESETn VGND VGND VPWR VPWR _23342_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18836__B1 _16518_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22632__B2 _22922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12258__A2_N _24761_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25188_ _24942_/CLK _25188_/D HRESETn VGND VGND VPWR VPWR _25188_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_123_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12153_ _12153_/A VGND VGND VPWR VPWR _12153_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12912__D _12903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24139_ _24136_/CLK _18725_/Y HRESETn VGND VGND VPWR VPWR _24139_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12084_ _12083_/Y _12079_/X _11853_/X _12079_/X VGND VGND VPWR VPWR _12084_/X sky130_fd_sc_hd__a2bb2o_4
X_16961_ _24709_/Q _16960_/Y _16007_/Y _24387_/Q VGND VGND VPWR VPWR _16961_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18700_ _18599_/X _18701_/B VGND VGND VPWR VPWR _18700_/X sky130_fd_sc_hd__or2_4
X_15912_ _24771_/Q _13540_/B VGND VGND VPWR VPWR _15912_/X sky130_fd_sc_hd__or2_4
X_19680_ _23645_/Q VGND VGND VPWR VPWR _19680_/Y sky130_fd_sc_hd__inv_2
X_16892_ _22181_/A VGND VGND VPWR VPWR _17867_/A sky130_fd_sc_hd__inv_2
XFILLER_42_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25235__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18631_ _18683_/A VGND VGND VPWR VPWR _18792_/A sky130_fd_sc_hd__buf_2
XANTENNA__17272__C1 _17271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15843_ _15843_/A _15703_/A VGND VGND VPWR VPWR _15843_/X sky130_fd_sc_hd__or2_4
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15822__B1 _24820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18562_ _18393_/Y _18562_/B VGND VGND VPWR VPWR _18575_/B sky130_fd_sc_hd__or2_4
X_12986_ _12299_/Y _13030_/A VGND VGND VPWR VPWR _12999_/C sky130_fd_sc_hd__or2_4
X_15774_ _15845_/A VGND VGND VPWR VPWR _15774_/X sky130_fd_sc_hd__buf_2
XFILLER_80_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17513_ _11831_/A _17512_/A _11831_/Y _17512_/Y VGND VGND VPWR VPWR _17513_/X sky130_fd_sc_hd__o22a_4
X_14725_ _25054_/Q VGND VGND VPWR VPWR _14725_/Y sky130_fd_sc_hd__inv_2
X_11937_ _11937_/A VGND VGND VPWR VPWR _19622_/A sky130_fd_sc_hd__buf_2
X_18493_ _18414_/A _18493_/B VGND VGND VPWR VPWR _18495_/B sky130_fd_sc_hd__or2_4
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14389__B1 _13840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11841__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17444_ _17438_/Y _17441_/Y _17443_/X _17441_/Y VGND VGND VPWR VPWR _17444_/X sky130_fd_sc_hd__a2bb2o_4
X_11868_ _11864_/Y _11741_/X _11867_/X _11741_/X VGND VGND VPWR VPWR _11868_/X sky130_fd_sc_hd__a2bb2o_4
X_14656_ _25061_/Q VGND VGND VPWR VPWR _14656_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24870__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13607_ _14785_/A _13605_/B _13606_/Y VGND VGND VPWR VPWR _13626_/B sky130_fd_sc_hd__o21a_4
X_17375_ _17374_/X VGND VGND VPWR VPWR _17375_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17327__B1 _17279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11799_ HWDATA[15] VGND VGND VPWR VPWR _11800_/A sky130_fd_sc_hd__buf_2
X_14587_ _25081_/Q _14571_/A VGND VGND VPWR VPWR _14587_/X sky130_fd_sc_hd__or2_4
XANTENNA__21123__B2 _21335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19114_ _23841_/Q VGND VGND VPWR VPWR _19114_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24188__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16326_ _16322_/Y _16324_/X _16325_/X _16324_/X VGND VGND VPWR VPWR _16326_/X sky130_fd_sc_hd__a2bb2o_4
X_13538_ _25289_/Q VGND VGND VPWR VPWR _14620_/D sky130_fd_sc_hd__inv_2
XFILLER_9_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21050__A _21024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24117__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19045_ _19052_/A VGND VGND VPWR VPWR _19045_/X sky130_fd_sc_hd__buf_2
X_13469_ _13468_/X VGND VGND VPWR VPWR _13533_/B sky130_fd_sc_hd__buf_2
X_16257_ _16256_/Y _16254_/X _16064_/X _16254_/X VGND VGND VPWR VPWR _24639_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15208_ _15246_/A VGND VGND VPWR VPWR _15216_/A sky130_fd_sc_hd__buf_2
XANTENNA__18827__B1 _16469_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16188_ _16179_/Y _16187_/X _11743_/X _16187_/X VGND VGND VPWR VPWR _16188_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15139_ _15374_/A VGND VGND VPWR VPWR _15139_/Y sky130_fd_sc_hd__inv_2
X_19947_ _23549_/Q VGND VGND VPWR VPWR _19947_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22387__B1 _13557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19878_ _21788_/B _19873_/X _19625_/X _19873_/X VGND VGND VPWR VPWR _19878_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12875__B1 _12874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18829_ _16476_/Y _18603_/X _16476_/Y _18603_/X VGND VGND VPWR VPWR _18833_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15813__B1 _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21840_ _14483_/Y _14258_/A VGND VGND VPWR VPWR _21840_/X sky130_fd_sc_hd__or2_4
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14962__A2_N _24416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24958__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21771_ _21624_/A _21769_/X _21770_/X VGND VGND VPWR VPWR _21771_/X sky130_fd_sc_hd__and3_4
XFILLER_64_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11751__A _11777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23510_ _25055_/CLK _23510_/D VGND VGND VPWR VPWR _23510_/Q sky130_fd_sc_hd__dfxtp_4
X_20722_ _13131_/B VGND VGND VPWR VPWR _20722_/Y sky130_fd_sc_hd__inv_2
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24490_ _24447_/CLK _16661_/X HRESETn VGND VGND VPWR VPWR _24490_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15041__B2 _24444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23441_ _23441_/CLK _23441_/D VGND VGND VPWR VPWR _20240_/A sky130_fd_sc_hd__dfxtp_4
X_20653_ _20652_/X VGND VGND VPWR VPWR _23979_/D sky130_fd_sc_hd__inv_2
Xclkbuf_7_100_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_201_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17318__B1 _17271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12285__C _12285_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24540__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23372_ _23904_/CLK _23372_/D VGND VGND VPWR VPWR _23372_/Q sky130_fd_sc_hd__dfxtp_4
X_20584_ _23942_/Q _18879_/X _20583_/Y _20556_/A VGND VGND VPWR VPWR _20584_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22056__A _22055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25111_ _23959_/CLK _14467_/X HRESETn VGND VGND VPWR VPWR _14465_/A sky130_fd_sc_hd__dfrtp_4
X_22323_ _22316_/Y _22318_/Y _22319_/X _22322_/Y _21547_/Y VGND VGND VPWR VPWR _22323_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_136_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25042_ _25043_/CLK _14830_/X HRESETn VGND VGND VPWR VPWR _25042_/Q sky130_fd_sc_hd__dfrtp_4
X_22254_ _21454_/A _22254_/B _22254_/C VGND VGND VPWR VPWR _22255_/C sky130_fd_sc_hd__and3_4
XANTENNA__15895__A3 _11818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21205_ _13780_/X _21203_/X _21162_/A _21204_/X VGND VGND VPWR VPWR _21205_/X sky130_fd_sc_hd__a211o_4
XFILLER_133_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22185_ _25513_/Q _22407_/B _21103_/A _22184_/X VGND VGND VPWR VPWR _22186_/C sky130_fd_sc_hd__a211o_4
X_21136_ _12123_/Y _21014_/A _12054_/A _21135_/Y VGND VGND VPWR VPWR _21137_/B sky130_fd_sc_hd__a211o_4
XANTENNA__20304__A _20298_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11926__A _11947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21067_ _21067_/A VGND VGND VPWR VPWR _21067_/X sky130_fd_sc_hd__buf_2
XFILLER_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21119__B _21333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20928__B2 _20913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20018_ _23525_/Q VGND VGND VPWR VPWR _20018_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15804__B1 _24833_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12840_ _25383_/Q VGND VGND VPWR VPWR _12840_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24826_ _24868_/CLK _24826_/D HRESETn VGND VGND VPWR VPWR _24826_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22145__A3 _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24699__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12771_ _12771_/A VGND VGND VPWR VPWR _12841_/B sky130_fd_sc_hd__inv_2
X_21969_ _21969_/A _21995_/A VGND VGND VPWR VPWR _21969_/X sky130_fd_sc_hd__or2_4
XANTENNA__21353__A1 _14876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24757_ _24759_/CLK _24757_/D HRESETn VGND VGND VPWR VPWR _24757_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _13787_/A _12057_/A VGND VGND VPWR VPWR _13813_/A sky130_fd_sc_hd__or2_4
X_14510_ _23952_/Q VGND VGND VPWR VPWR _14510_/X sky130_fd_sc_hd__buf_2
XANTENNA__24628__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15516_/A VGND VGND VPWR VPWR _15490_/X sky130_fd_sc_hd__buf_2
X_23708_ _23683_/CLK _23708_/D VGND VGND VPWR VPWR _23708_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24688_ _24692_/CLK _24688_/D HRESETn VGND VGND VPWR VPWR _16115_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15032__B2 _15023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11653_/A VGND VGND VPWR VPWR _11701_/A sky130_fd_sc_hd__inv_2
X_14441_ _25122_/Q VGND VGND VPWR VPWR _14441_/Y sky130_fd_sc_hd__inv_2
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23639_ _24288_/CLK _23639_/D VGND VGND VPWR VPWR _19696_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24281__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14372_ _25141_/Q _14330_/X _14356_/X _12090_/A _14354_/Y VGND VGND VPWR VPWR _14372_/X
+ sky130_fd_sc_hd__a32o_4
X_17160_ _17160_/A _17160_/B _17160_/C VGND VGND VPWR VPWR _17160_/X sky130_fd_sc_hd__and3_4
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13323_ _13162_/A VGND VGND VPWR VPWR _13461_/A sky130_fd_sc_hd__buf_2
X_16111_ _16110_/Y _16106_/X _15952_/X _16106_/X VGND VGND VPWR VPWR _16111_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25309_ _25309_/CLK _25309_/D HRESETn VGND VGND VPWR VPWR _13481_/A sky130_fd_sc_hd__dfrtp_4
X_17091_ _17023_/Y _17091_/B VGND VGND VPWR VPWR _17091_/X sky130_fd_sc_hd__or2_4
XFILLER_52_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12197__A2_N _24735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13254_ _13168_/A _13254_/B _13253_/X VGND VGND VPWR VPWR _13254_/X sky130_fd_sc_hd__and3_4
X_16042_ _16042_/A VGND VGND VPWR VPWR _16042_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25487__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12205_ _12202_/A _24743_/Q _12203_/X _12204_/Y VGND VGND VPWR VPWR _12212_/B sky130_fd_sc_hd__o22a_4
XANTENNA__20616__B1 _20662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13185_ _13181_/X _13184_/X _13162_/X VGND VGND VPWR VPWR _13185_/X sky130_fd_sc_hd__o21a_4
XFILLER_135_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25416__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19801_ _13171_/B VGND VGND VPWR VPWR _19801_/Y sky130_fd_sc_hd__inv_2
X_12136_ _12116_/A _12125_/A _12116_/A _12125_/A VGND VGND VPWR VPWR _12136_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17993_ _18224_/A _17993_/B _17993_/C VGND VGND VPWR VPWR _17994_/C sky130_fd_sc_hd__or3_4
X_19732_ _23627_/Q VGND VGND VPWR VPWR _19732_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12067_ _12057_/A VGND VGND VPWR VPWR _13789_/B sky130_fd_sc_hd__buf_2
X_16944_ _24690_/Q _16943_/Y _16115_/Y _16941_/A VGND VGND VPWR VPWR _16944_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16048__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21041__B1 _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19663_ _19676_/A VGND VGND VPWR VPWR _19663_/X sky130_fd_sc_hd__buf_2
X_16875_ _19790_/A VGND VGND VPWR VPWR _16875_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18619__A _24121_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18614_ _18679_/A VGND VGND VPWR VPWR _18614_/X sky130_fd_sc_hd__buf_2
XFILLER_64_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_129_0_HCLK clkbuf_7_64_0_HCLK/X VGND VGND VPWR VPWR _23887_/CLK sky130_fd_sc_hd__clkbuf_1
X_15826_ _15829_/A VGND VGND VPWR VPWR _15826_/X sky130_fd_sc_hd__buf_2
X_19594_ _22046_/A _19588_/X _19407_/X _19593_/X VGND VGND VPWR VPWR _23674_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18545_ _24160_/Q _18545_/B VGND VGND VPWR VPWR _18546_/C sky130_fd_sc_hd__or2_4
XFILLER_52_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15757_ _12549_/Y _15754_/X _15756_/X _15754_/X VGND VGND VPWR VPWR _15757_/X sky130_fd_sc_hd__a2bb2o_4
X_12969_ _12969_/A VGND VGND VPWR VPWR _25359_/D sky130_fd_sc_hd__inv_2
XANTENNA__17548__B1 _11844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21344__A1 SSn_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22541__B1 _22527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24369__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14708_ _14707_/Y VGND VGND VPWR VPWR _14708_/X sky130_fd_sc_hd__buf_2
XFILLER_61_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18476_ _18476_/A _18476_/B _18476_/C VGND VGND VPWR VPWR _18477_/C sky130_fd_sc_hd__or3_4
X_15688_ _15677_/X _15684_/A _14620_/B _15682_/C _15687_/X VGND VGND VPWR VPWR _15689_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16220__B1 _15962_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17427_ _24317_/Q VGND VGND VPWR VPWR _17427_/Y sky130_fd_sc_hd__inv_2
X_14639_ _14785_/A VGND VGND VPWR VPWR _18202_/A sky130_fd_sc_hd__buf_2
XFILLER_127_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17358_ _17350_/B _17349_/X VGND VGND VPWR VPWR _17361_/B sky130_fd_sc_hd__or2_4
X_16309_ _16308_/Y _16303_/X _15952_/X _16303_/X VGND VGND VPWR VPWR _16309_/X sky130_fd_sc_hd__a2bb2o_4
X_17289_ _17289_/A _17284_/B _17288_/X VGND VGND VPWR VPWR _17289_/X sky130_fd_sc_hd__or3_4
X_19028_ _19027_/Y _19023_/X _18977_/X _19023_/X VGND VGND VPWR VPWR _19028_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15877__A3 _15729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20607__B1 _20662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23933__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23138__C _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11746__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19225__B1 _19133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13664__C _20900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23990_ _23989_/CLK _20671_/X HRESETn VGND VGND VPWR VPWR _23990_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16561__A1_N _16560_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_25_0_HCLK clkbuf_7_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22941_ _24723_/Q _21021_/X _21050_/X _22940_/X VGND VGND VPWR VPWR _22941_/X sky130_fd_sc_hd__a211o_4
XFILLER_99_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_88_0_HCLK clkbuf_6_44_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_88_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22872_ _22872_/A _22872_/B VGND VGND VPWR VPWR _22872_/X sky130_fd_sc_hd__and2_4
X_21823_ _21707_/X _21744_/X _21784_/X _21822_/X VGND VGND VPWR VPWR HRDATA[3] sky130_fd_sc_hd__or4_4
XFILLER_83_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24792__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24611_ _24885_/CLK _16335_/X HRESETn VGND VGND VPWR VPWR _24611_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16049__A _24713_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24721__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24542_ _24541_/CLK _24542_/D HRESETn VGND VGND VPWR VPWR _16518_/A sky130_fd_sc_hd__dfrtp_4
X_21754_ _21609_/A _21752_/X _21753_/X VGND VGND VPWR VPWR _21754_/X sky130_fd_sc_hd__and3_4
XFILLER_70_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24039__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20705_ _20704_/X VGND VGND VPWR VPWR _20705_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23170__A _23170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24473_ _24581_/CLK _24473_/D HRESETn VGND VGND VPWR VPWR _24473_/Q sky130_fd_sc_hd__dfrtp_4
X_21685_ _21495_/X _21684_/X _11694_/Y _21495_/X VGND VGND VPWR VPWR _21685_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23424_ _24923_/CLK _20286_/X VGND VGND VPWR VPWR _20285_/A sky130_fd_sc_hd__dfxtp_4
X_20636_ _14241_/Y _20628_/X _20619_/X _20635_/X VGND VGND VPWR VPWR _20637_/A sky130_fd_sc_hd__a211o_4
XFILLER_138_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23355_ _23342_/X VGND VGND VPWR VPWR IRQ[1] sky130_fd_sc_hd__buf_2
X_20567_ _18876_/X _20567_/B _20571_/C VGND VGND VPWR VPWR _20567_/X sky130_fd_sc_hd__and3_4
XANTENNA__15317__A2 _15316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22306_ _22306_/A VGND VGND VPWR VPWR _22306_/Y sky130_fd_sc_hd__inv_2
X_23286_ _15559_/Y _22872_/B VGND VGND VPWR VPWR _23286_/X sky130_fd_sc_hd__and2_4
X_20498_ _23995_/Q _20512_/B _20497_/X VGND VGND VPWR VPWR _20498_/X sky130_fd_sc_hd__a21o_4
X_25025_ _25024_/CLK _25025_/D HRESETn VGND VGND VPWR VPWR _25025_/Q sky130_fd_sc_hd__dfrtp_4
X_22237_ _22229_/A _19892_/Y VGND VGND VPWR VPWR _22237_/X sky130_fd_sc_hd__or2_4
XFILLER_133_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21271__B1 _21270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22168_ _13503_/Y _12097_/X _12031_/Y _12071_/A VGND VGND VPWR VPWR _22168_/X sky130_fd_sc_hd__o22a_4
XFILLER_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21119_ _21119_/A _21333_/A VGND VGND VPWR VPWR _21119_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__23012__A1 _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14990_ _14990_/A VGND VGND VPWR VPWR _15283_/A sky130_fd_sc_hd__inv_2
X_22099_ _22098_/X VGND VGND VPWR VPWR _22101_/C sky130_fd_sc_hd__inv_2
XFILLER_130_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13941_ _13889_/C VGND VGND VPWR VPWR _13941_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13871__A _23989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24809__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16660_ _24490_/Q VGND VGND VPWR VPWR _16660_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13872_ _22111_/A _13861_/X _21829_/A _13863_/X VGND VGND VPWR VPWR _13872_/X sky130_fd_sc_hd__o22a_4
XFILLER_47_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15611_ _15611_/A VGND VGND VPWR VPWR _22559_/A sky130_fd_sc_hd__inv_2
XANTENNA__19519__B2 _19516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12823_ _12854_/A _24798_/Q _25375_/Q _12822_/Y VGND VGND VPWR VPWR _12823_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13590__B _14555_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24809_ _24836_/CLK _24809_/D HRESETn VGND VGND VPWR VPWR _24809_/Q sky130_fd_sc_hd__dfrtp_4
X_16591_ _16590_/Y _16588_/X _16235_/X _16588_/X VGND VGND VPWR VPWR _24515_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12487__A _12278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18330_ _19105_/A _18326_/X _18329_/X VGND VGND VPWR VPWR _18330_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__24462__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15542_ _15542_/A VGND VGND VPWR VPWR _15542_/Y sky130_fd_sc_hd__inv_2
X_12754_ _12753_/X _24788_/Q _12753_/X _24788_/Q VGND VGND VPWR VPWR _12754_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11705_ _11647_/X _11652_/X _17445_/C _11967_/C VGND VGND VPWR VPWR _11705_/X sky130_fd_sc_hd__o22a_4
X_18261_ _18261_/A _18230_/B VGND VGND VPWR VPWR _18262_/A sky130_fd_sc_hd__or2_4
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12679_/A _12689_/B VGND VGND VPWR VPWR _12685_/Y sky130_fd_sc_hd__nand2_4
X_15473_ _24941_/Q VGND VGND VPWR VPWR _15473_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23079__B2 _22827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _16332_/Y _17248_/A _16332_/Y _17248_/A VGND VGND VPWR VPWR _17212_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14424_ _14423_/Y _14419_/X _14403_/X _14419_/X VGND VGND VPWR VPWR _25128_/D sky130_fd_sc_hd__a2bb2o_4
X_18192_ _18058_/A _18192_/B _18192_/C VGND VGND VPWR VPWR _18192_/X sky130_fd_sc_hd__or3_4
XFILLER_128_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20209__A _20209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17143_ _17143_/A _17134_/B _17143_/C VGND VGND VPWR VPWR _17143_/X sky130_fd_sc_hd__and3_4
XANTENNA__22127__C _22127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14355_ _14354_/Y VGND VGND VPWR VPWR _14355_/X sky130_fd_sc_hd__buf_2
XFILLER_128_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15310__B _15310_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13306_ _13454_/A _13300_/X _13305_/X VGND VGND VPWR VPWR _13306_/X sky130_fd_sc_hd__or3_4
X_14286_ _25170_/Q _13643_/B VGND VGND VPWR VPWR _25170_/D sky130_fd_sc_hd__and2_4
X_17074_ _17066_/B _17065_/X _17026_/Y VGND VGND VPWR VPWR _17075_/C sky130_fd_sc_hd__o21a_4
X_13237_ _13317_/A _13237_/B VGND VGND VPWR VPWR _13238_/C sky130_fd_sc_hd__or2_4
X_16025_ _16024_/Y _16022_/X _15957_/X _16022_/X VGND VGND VPWR VPWR _16025_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23251__A1 _12385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19455__B1 _19364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25250__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16269__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15738__A1_N _12559_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13168_ _13168_/A VGND VGND VPWR VPWR _13191_/A sky130_fd_sc_hd__buf_2
XFILLER_3_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12119_ _12119_/A VGND VGND VPWR VPWR _12119_/X sky130_fd_sc_hd__buf_2
XANTENNA__19207__B1 _19206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13099_ _13042_/A VGND VGND VPWR VPWR _13115_/C sky130_fd_sc_hd__buf_2
X_17976_ _17990_/A VGND VGND VPWR VPWR _18104_/A sky130_fd_sc_hd__buf_2
XFILLER_85_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19715_ _15766_/A VGND VGND VPWR VPWR _19715_/X sky130_fd_sc_hd__buf_2
X_16927_ _16927_/A VGND VGND VPWR VPWR _16927_/X sky130_fd_sc_hd__buf_2
XFILLER_133_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22762__B1 _24823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19646_ _19638_/Y VGND VGND VPWR VPWR _19646_/X sky130_fd_sc_hd__buf_2
X_16858_ _19777_/A VGND VGND VPWR VPWR _16858_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15809_ _15809_/A VGND VGND VPWR VPWR _15809_/X sky130_fd_sc_hd__buf_2
X_19577_ _19576_/Y _19574_/X _11955_/X _19574_/X VGND VGND VPWR VPWR _23678_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16789_ _15010_/Y _16783_/X _16442_/X _16783_/X VGND VGND VPWR VPWR _16789_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12397__A _12385_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22514__B1 _21106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18528_ _18541_/A _18526_/X _18527_/X VGND VGND VPWR VPWR _24166_/D sky130_fd_sc_hd__and3_4
XANTENNA__21868__A2 _21418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24132__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18459_ _18459_/A VGND VGND VPWR VPWR _18460_/A sky130_fd_sc_hd__inv_2
XFILLER_107_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18084__A _18046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21470_ _17706_/A VGND VGND VPWR VPWR _21649_/A sky130_fd_sc_hd__buf_2
XANTENNA__22817__A1 _24720_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20421_ _20421_/A VGND VGND VPWR VPWR _23920_/D sky130_fd_sc_hd__buf_2
XFILLER_88_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12230__B2 _22141_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25338__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23140_ _24761_/Q _23140_/B VGND VGND VPWR VPWR _23140_/X sky130_fd_sc_hd__or2_4
X_20352_ _20339_/Y VGND VGND VPWR VPWR _20352_/X sky130_fd_sc_hd__buf_2
XFILLER_106_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23071_ _22808_/X _23071_/B _23071_/C VGND VGND VPWR VPWR _23071_/X sky130_fd_sc_hd__and3_4
X_20283_ _20290_/A VGND VGND VPWR VPWR _20283_/X sky130_fd_sc_hd__buf_2
XFILLER_115_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16332__A _24612_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22022_ _21671_/A _22022_/B _22021_/X VGND VGND VPWR VPWR _22022_/X sky130_fd_sc_hd__and3_4
XFILLER_66_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24973__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13494__B1 _13472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23973_ _24943_/CLK _20627_/Y HRESETn VGND VGND VPWR VPWR _23973_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14787__A _18177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24902__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22924_ _16490_/A _22879_/X _22798_/X VGND VGND VPWR VPWR _22924_/X sky130_fd_sc_hd__o21a_4
XFILLER_60_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16432__B1 _16057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_112_0_HCLK clkbuf_7_56_0_HCLK/X VGND VGND VPWR VPWR _24159_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21308__A1 _21275_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22855_ _22759_/X _22853_/X _22854_/X _24825_/Q _22761_/X VGND VGND VPWR VPWR _22856_/B
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_8_175_0_HCLK clkbuf_7_87_0_HCLK/X VGND VGND VPWR VPWR _23711_/CLK sky130_fd_sc_hd__clkbuf_1
X_21806_ _21802_/X _21805_/X _21481_/X VGND VGND VPWR VPWR _21806_/X sky130_fd_sc_hd__o21a_4
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22786_ _22786_/A VGND VGND VPWR VPWR _22786_/X sky130_fd_sc_hd__buf_2
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21737_ _21731_/X _21737_/B VGND VGND VPWR VPWR _21737_/Y sky130_fd_sc_hd__nor2_4
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24525_ _24557_/CLK _24525_/D HRESETn VGND VGND VPWR VPWR _24525_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23331__C _23331_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12470_ _12278_/C _12469_/X VGND VGND VPWR VPWR _12471_/D sky130_fd_sc_hd__or2_4
X_21668_ _21668_/A VGND VGND VPWR VPWR _21671_/A sky130_fd_sc_hd__buf_2
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24456_ _24457_/CLK _24456_/D HRESETn VGND VGND VPWR VPWR _16745_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20029__A _20036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20619_ _20619_/A VGND VGND VPWR VPWR _20619_/X sky130_fd_sc_hd__buf_2
X_23407_ _24209_/CLK _23407_/D VGND VGND VPWR VPWR _20329_/A sky130_fd_sc_hd__dfxtp_4
X_24387_ _24391_/CLK _17073_/X HRESETn VGND VGND VPWR VPWR _24387_/Q sky130_fd_sc_hd__dfrtp_4
X_21599_ _21631_/A _21599_/B _21599_/C VGND VGND VPWR VPWR _21599_/X sky130_fd_sc_hd__and3_4
XANTENNA__15537__A2_N _15535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25079__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14140_ _14139_/X VGND VGND VPWR VPWR _14140_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23985__D sda_i_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23338_ _25258_/Q _23337_/X VGND VGND VPWR VPWR _23338_/X sky130_fd_sc_hd__and2_4
XANTENNA__19537__B _16725_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25008__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14071_ _14054_/Y _14071_/B _14050_/X _14015_/X VGND VGND VPWR VPWR _14071_/X sky130_fd_sc_hd__or4_4
XFILLER_125_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23269_ _24765_/Q _23269_/B VGND VGND VPWR VPWR _23269_/X sky130_fd_sc_hd__or2_4
XFILLER_106_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16242__A _11818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13022_ _25349_/Q _13026_/B VGND VGND VPWR VPWR _13024_/B sky130_fd_sc_hd__or2_4
X_25008_ _25010_/CLK _25008_/D HRESETn VGND VGND VPWR VPWR _15241_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_121_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17830_ _17755_/Y _17830_/B VGND VGND VPWR VPWR _17833_/B sky130_fd_sc_hd__or2_4
XANTENNA__19553__A _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17761_ _17741_/Y _16943_/Y _17761_/C _17792_/B VGND VGND VPWR VPWR _17761_/X sky130_fd_sc_hd__or4_4
X_14973_ _25017_/Q _14971_/Y _15212_/A _14969_/A VGND VGND VPWR VPWR _14973_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13485__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19500_ _19494_/Y VGND VGND VPWR VPWR _19500_/X sky130_fd_sc_hd__buf_2
XANTENNA__22744__B1 _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16712_ _16645_/A VGND VGND VPWR VPWR _16712_/X sky130_fd_sc_hd__buf_2
XANTENNA__24643__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13924_ _13924_/A VGND VGND VPWR VPWR _13924_/X sky130_fd_sc_hd__buf_2
X_17692_ _17692_/A _17691_/X _17681_/X VGND VGND VPWR VPWR _17692_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_71_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_71_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19431_ _19431_/A VGND VGND VPWR VPWR _19431_/X sky130_fd_sc_hd__buf_2
X_16643_ _16643_/A VGND VGND VPWR VPWR _16643_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13855_ _13850_/Y VGND VGND VPWR VPWR _13855_/X sky130_fd_sc_hd__buf_2
XFILLER_63_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12806_ _12806_/A VGND VGND VPWR VPWR _22660_/A sky130_fd_sc_hd__buf_2
X_19362_ _19360_/Y _19356_/X _19294_/X _19361_/X VGND VGND VPWR VPWR _19362_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12105__A1_N _12104_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16574_ _24521_/Q VGND VGND VPWR VPWR _16574_/Y sky130_fd_sc_hd__inv_2
X_13786_ _13786_/A VGND VGND VPWR VPWR _23336_/A sky130_fd_sc_hd__inv_2
X_18313_ _17729_/Y _24202_/Q _17729_/A _21196_/A VGND VGND VPWR VPWR _18314_/A sky130_fd_sc_hd__o22a_4
XFILLER_128_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15525_ _15523_/Y _15524_/X HADDR[9] _15524_/X VGND VGND VPWR VPWR _24921_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12737_ _12737_/A _12736_/X _12721_/X VGND VGND VPWR VPWR _25389_/D sky130_fd_sc_hd__and3_4
X_19293_ _13282_/B VGND VGND VPWR VPWR _19293_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18244_ _22532_/A _18242_/X _11821_/X _18242_/X VGND VGND VPWR VPWR _24223_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21305__A2_N _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15456_ _14279_/A VGND VGND VPWR VPWR _20602_/A sky130_fd_sc_hd__buf_2
X_12668_ _12670_/B VGND VGND VPWR VPWR _12669_/B sky130_fd_sc_hd__inv_2
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _14407_/A VGND VGND VPWR VPWR _14475_/B sky130_fd_sc_hd__buf_2
X_18175_ _18175_/A _18982_/A VGND VGND VPWR VPWR _18176_/C sky130_fd_sc_hd__or2_4
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22275__A2 _22269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15387_ _15092_/Y _15387_/B VGND VGND VPWR VPWR _15421_/A sky130_fd_sc_hd__or2_4
X_12599_ _12569_/X _12599_/B _12599_/C _12598_/X VGND VGND VPWR VPWR _12600_/B sky130_fd_sc_hd__or4_4
XANTENNA__25431__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17126_ _17126_/A VGND VGND VPWR VPWR _24372_/D sky130_fd_sc_hd__inv_2
XFILLER_117_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14338_ _14338_/A VGND VGND VPWR VPWR _14338_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22680__C1 _22675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17057_ _17022_/Y _17051_/B _17053_/B _17056_/X VGND VGND VPWR VPWR _17057_/X sky130_fd_sc_hd__a211o_4
X_14269_ _14268_/Y _14264_/X _13800_/X _14264_/X VGND VGND VPWR VPWR _14269_/X sky130_fd_sc_hd__a2bb2o_4
X_16008_ _16007_/Y _16003_/X _15944_/X _16003_/X VGND VGND VPWR VPWR _16008_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21993__A _13784_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17959_ _18059_/A _17951_/X _17958_/X _15677_/X _15685_/X VGND VGND VPWR VPWR _17959_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_97_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24384__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20970_ scl_oen_o_S4 _20970_/B VGND VGND VPWR VPWR _20970_/X sky130_fd_sc_hd__and2_4
XANTENNA__19600__B1 _19599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24313__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19629_ _19629_/A VGND VGND VPWR VPWR _19629_/X sky130_fd_sc_hd__buf_2
XFILLER_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22640_ _12799_/X _22565_/X _22639_/X VGND VGND VPWR VPWR _22640_/X sky130_fd_sc_hd__o21a_4
XFILLER_0_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_248_0_HCLK clkbuf_7_124_0_HCLK/X VGND VGND VPWR VPWR _24852_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22329__A _21942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22571_ _24578_/Q _22522_/B VGND VGND VPWR VPWR _22571_/X sky130_fd_sc_hd__or2_4
XFILLER_90_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25519__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21522_ _23306_/A _21521_/X VGND VGND VPWR VPWR _21522_/X sky130_fd_sc_hd__and2_4
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24310_ _24208_/CLK _24310_/D HRESETn VGND VGND VPWR VPWR _24310_/Q sky130_fd_sc_hd__dfrtp_4
X_25290_ _25290_/CLK _13537_/X HRESETn VGND VGND VPWR VPWR _13536_/A sky130_fd_sc_hd__dfrtp_4
X_24241_ _24186_/CLK _17910_/X HRESETn VGND VGND VPWR VPWR _17909_/A sky130_fd_sc_hd__dfrtp_4
X_21453_ _21191_/A VGND VGND VPWR VPWR _21454_/A sky130_fd_sc_hd__buf_2
XFILLER_21_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25172__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20404_ _23376_/Q VGND VGND VPWR VPWR _20404_/Y sky130_fd_sc_hd__inv_2
X_24172_ _24502_/CLK _18504_/X HRESETn VGND VGND VPWR VPWR _24172_/Q sky130_fd_sc_hd__dfrtp_4
X_21384_ _21381_/A _21384_/B VGND VGND VPWR VPWR _21384_/X sky130_fd_sc_hd__or2_4
XANTENNA__25101__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23123_ _23119_/X _23120_/X _23121_/X _23122_/X VGND VGND VPWR VPWR _23124_/B sky130_fd_sc_hd__o22a_4
X_20335_ _20335_/A VGND VGND VPWR VPWR _20335_/Y sky130_fd_sc_hd__inv_2
X_23054_ _23054_/A _23053_/X VGND VGND VPWR VPWR _23054_/Y sky130_fd_sc_hd__nor2_4
X_20266_ _20266_/A VGND VGND VPWR VPWR _20266_/X sky130_fd_sc_hd__buf_2
XANTENNA__21777__A1 _21759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22005_ _22009_/A VGND VGND VPWR VPWR _22005_/X sky130_fd_sc_hd__buf_2
XFILLER_62_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20197_ _20195_/Y _20191_/X _16872_/A _20196_/X VGND VGND VPWR VPWR _23458_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21408__A _21408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11970_ _11958_/X _17445_/C _11970_/C _11970_/D VGND VGND VPWR VPWR _11970_/X sky130_fd_sc_hd__or4_4
X_23956_ _23989_/CLK _23956_/D HRESETn VGND VGND VPWR VPWR _23956_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24054__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_58_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22907_ _12286_/C _22489_/X _24264_/Q _22906_/X VGND VGND VPWR VPWR _22907_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12690__A1 _12567_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23887_ _23887_/CLK _18981_/X VGND VGND VPWR VPWR _18980_/A sky130_fd_sc_hd__dfxtp_4
X_13640_ _13526_/Y VGND VGND VPWR VPWR _13640_/X sky130_fd_sc_hd__buf_2
XFILLER_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22838_ _23021_/A _22832_/X _22838_/C VGND VGND VPWR VPWR _22838_/X sky130_fd_sc_hd__and3_4
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21143__A _21143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _25255_/Q _13568_/X _13569_/Y _13570_/Y VGND VGND VPWR VPWR _13578_/B sky130_fd_sc_hd__o22a_4
XFILLER_72_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12442__A1 _12286_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22769_ _22419_/X VGND VGND VPWR VPWR _22769_/X sky130_fd_sc_hd__buf_2
X_15310_ _15155_/Y _15310_/B _15309_/X VGND VGND VPWR VPWR _15313_/B sky130_fd_sc_hd__or3_4
XFILLER_34_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _12679_/A _24858_/Q _12520_/Y _24858_/Q VGND VGND VPWR VPWR _12531_/A sky130_fd_sc_hd__a2bb2o_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24508_ _24120_/CLK _24508_/D HRESETn VGND VGND VPWR VPWR _16608_/A sky130_fd_sc_hd__dfrtp_4
X_16290_ _16287_/Y _16282_/X _15940_/X _16289_/X VGND VGND VPWR VPWR _16290_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25488_ _25488_/CLK _11968_/X HRESETn VGND VGND VPWR VPWR _11961_/A sky130_fd_sc_hd__dfrtp_4
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15241_ _15241_/A _15240_/Y VGND VGND VPWR VPWR _15243_/B sky130_fd_sc_hd__or2_4
X_12453_ _12455_/B VGND VGND VPWR VPWR _12454_/B sky130_fd_sc_hd__inv_2
XFILLER_138_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24439_ _24407_/CLK _16779_/X HRESETn VGND VGND VPWR VPWR _24439_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18452__A _18743_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12384_ _12391_/A _13008_/B VGND VGND VPWR VPWR _12397_/B sky130_fd_sc_hd__or2_4
X_15172_ _15165_/A _15171_/X VGND VGND VPWR VPWR _15172_/X sky130_fd_sc_hd__or2_4
X_14123_ _14181_/B _14129_/A VGND VGND VPWR VPWR _14124_/A sky130_fd_sc_hd__and2_4
XFILLER_114_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19980_ _23538_/Q VGND VGND VPWR VPWR _22029_/B sky130_fd_sc_hd__inv_2
XFILLER_126_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18931_ _18929_/Y _18925_/X _17424_/X _18930_/X VGND VGND VPWR VPWR _23906_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24895__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14054_ _14053_/X VGND VGND VPWR VPWR _14054_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13005_ _12294_/Y _13005_/B VGND VGND VPWR VPWR _13005_/X sky130_fd_sc_hd__or2_4
XANTENNA__24824__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18862_ _16473_/Y _24139_/Q _16488_/Y _24133_/Q VGND VGND VPWR VPWR _18864_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19830__B1 _19783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16700__A _16645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17813_ _16900_/A _17813_/B VGND VGND VPWR VPWR _17815_/B sky130_fd_sc_hd__or2_4
X_18793_ _18608_/X _18792_/X _18724_/A _18788_/Y VGND VGND VPWR VPWR _18794_/A sky130_fd_sc_hd__a211o_4
XFILLER_130_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17744_ _17744_/A VGND VGND VPWR VPWR _17744_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15316__A _15310_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14956_ _14955_/Y VGND VGND VPWR VPWR _15193_/A sky130_fd_sc_hd__buf_2
XFILLER_94_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14220__A _14220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18397__B1 _16223_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13907_ _13906_/X VGND VGND VPWR VPWR _13908_/B sky130_fd_sc_hd__inv_2
X_17675_ _17652_/X _17672_/B _17675_/C VGND VGND VPWR VPWR _17675_/X sky130_fd_sc_hd__and3_4
X_14887_ _14886_/X _24412_/Q _14886_/X _24412_/Q VGND VGND VPWR VPWR _14887_/X sky130_fd_sc_hd__a2bb2o_4
X_19414_ _18139_/B VGND VGND VPWR VPWR _19414_/Y sky130_fd_sc_hd__inv_2
X_16626_ RsRx_S0 _16172_/B _16625_/Y VGND VGND VPWR VPWR _16634_/B sky130_fd_sc_hd__o21a_4
X_13838_ _13551_/Y _13833_/X _13837_/X _13833_/X VGND VGND VPWR VPWR _13838_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22149__A _22035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23142__B1 _24833_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19345_ _18150_/B VGND VGND VPWR VPWR _19345_/Y sky130_fd_sc_hd__inv_2
X_16557_ _24528_/Q VGND VGND VPWR VPWR _16557_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_1_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_13769_ _25263_/Q VGND VGND VPWR VPWR _13769_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22496__A2 _22442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16147__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_15_0_HCLK clkbuf_7_7_0_HCLK/X VGND VGND VPWR VPWR _24089_/CLK sky130_fd_sc_hd__clkbuf_1
X_15508_ _11729_/C VGND VGND VPWR VPWR _15508_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19276_ _21752_/B _19271_/X _16881_/X _19271_/X VGND VGND VPWR VPWR _23784_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16488_ _24554_/Q VGND VGND VPWR VPWR _16488_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_78_0_HCLK clkbuf_8_79_0_HCLK/A VGND VGND VPWR VPWR _25192_/CLK sky130_fd_sc_hd__clkbuf_1
X_18227_ _17960_/X _18226_/X _24229_/Q _18021_/A VGND VGND VPWR VPWR _24229_/D sky130_fd_sc_hd__o22a_4
X_15439_ _13924_/X _15437_/X _15432_/X _24961_/Q _15438_/X VGND VGND VPWR VPWR _15439_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15986__A _15986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19649__B1 _19547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18158_ _18056_/A _19210_/A VGND VGND VPWR VPWR _18158_/X sky130_fd_sc_hd__or2_4
X_17109_ _17034_/B _17105_/X VGND VGND VPWR VPWR _17109_/Y sky130_fd_sc_hd__nand2_4
XFILLER_116_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18089_ _18186_/A _19139_/A VGND VGND VPWR VPWR _18089_/X sky130_fd_sc_hd__or2_4
XFILLER_117_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20120_ _23486_/Q VGND VGND VPWR VPWR _21385_/B sky130_fd_sc_hd__inv_2
XFILLER_89_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22956__B1 _12584_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24565__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20051_ _22068_/B _20045_/X _19783_/X _20050_/X VGND VGND VPWR VPWR _23514_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18624__A1 _24509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17706__A _17706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11754__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23810_ _23818_/CLK _19204_/X VGND VGND VPWR VPWR _18056_/B sky130_fd_sc_hd__dfxtp_4
X_24790_ _24800_/CLK _15884_/X HRESETn VGND VGND VPWR VPWR _22857_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18388__B1 _24178_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20953_ _11991_/A _20953_/B VGND VGND VPWR VPWR _24085_/D sky130_fd_sc_hd__nor2_4
XFILLER_54_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23741_ _23446_/CLK _19397_/X VGND VGND VPWR VPWR _23741_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16938__B2 _16898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17441__A _14223_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _20889_/B VGND VGND VPWR VPWR _20884_/Y sky130_fd_sc_hd__inv_2
XPHY_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23672_ _23689_/CLK _23672_/D VGND VGND VPWR VPWR _19597_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22059__A _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25411_ _25411_/CLK _12660_/X HRESETn VGND VGND VPWR VPWR _12659_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22623_ _22623_/A _22587_/B VGND VGND VPWR VPWR _22623_/X sky130_fd_sc_hd__or2_4
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16057__A _16057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25353__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22554_ _21700_/X _22553_/X _21532_/X _24713_/Q _21299_/X VGND VGND VPWR VPWR _22554_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21695__B1 _24845_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25342_ _24852_/CLK _25342_/D HRESETn VGND VGND VPWR VPWR _25342_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17363__A1 _17350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21505_ _18272_/A _21500_/X _21502_/X _21504_/X VGND VGND VPWR VPWR _21505_/X sky130_fd_sc_hd__a211o_4
X_22485_ _21427_/X VGND VGND VPWR VPWR _22485_/X sky130_fd_sc_hd__buf_2
X_25273_ _25508_/CLK _13724_/X HRESETn VGND VGND VPWR VPWR _25273_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18272__A _18272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21436_ _23314_/B _21429_/X _23271_/A _21435_/X VGND VGND VPWR VPWR _21436_/Y sky130_fd_sc_hd__a22oi_4
X_24224_ _24346_/CLK _24224_/D HRESETn VGND VGND VPWR VPWR _24224_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17503__A2_N _17630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24155_ _24151_/CLK _18570_/X HRESETn VGND VGND VPWR VPWR _24155_/Q sky130_fd_sc_hd__dfrtp_4
X_21367_ _21264_/X _21363_/X _21365_/Y _21366_/X VGND VGND VPWR VPWR _21367_/X sky130_fd_sc_hd__a211o_4
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20318_ _19582_/X VGND VGND VPWR VPWR _20318_/X sky130_fd_sc_hd__buf_2
X_23106_ _21511_/X VGND VGND VPWR VPWR _23106_/X sky130_fd_sc_hd__buf_2
X_24086_ _25301_/CLK _20954_/X HRESETn VGND VGND VPWR VPWR _11991_/B sky130_fd_sc_hd__dfrtp_4
X_21298_ _22747_/B VGND VGND VPWR VPWR _23097_/A sky130_fd_sc_hd__buf_2
XFILLER_116_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23037_ _23034_/X _23036_/X _22968_/X _24865_/Q _22766_/X VGND VGND VPWR VPWR _23037_/X
+ sky130_fd_sc_hd__a32o_4
X_20249_ _23437_/Q VGND VGND VPWR VPWR _20249_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16520__A _24541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24235__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14810_ _14810_/A VGND VGND VPWR VPWR _14810_/X sky130_fd_sc_hd__buf_2
XFILLER_92_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15790_ _21025_/A VGND VGND VPWR VPWR _15791_/A sky130_fd_sc_hd__buf_2
XANTENNA__16641__A3 HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24988_ _24995_/CLK _24988_/D HRESETn VGND VGND VPWR VPWR _15080_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12112__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14741_ _14722_/X _14729_/Y _14740_/X _22036_/A _14723_/Y VGND VGND VPWR VPWR _25053_/D
+ sky130_fd_sc_hd__a32o_4
X_11953_ _11951_/Y _11947_/X _11952_/X _11947_/X VGND VGND VPWR VPWR _25491_/D sky130_fd_sc_hd__a2bb2o_4
X_23939_ _25122_/CLK _23939_/D HRESETn VGND VGND VPWR VPWR _23939_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21337__A1_N _14177_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25120__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17460_ _17459_/X _18344_/A _17459_/X _18344_/A VGND VGND VPWR VPWR _17489_/A sky130_fd_sc_hd__a2bb2o_4
X_14672_ _19152_/A _14671_/X _19152_/A _14671_/X VGND VGND VPWR VPWR _14672_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23072__B _21017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25183__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11884_ _11883_/Y _11878_/B VGND VGND VPWR VPWR _11884_/X sky130_fd_sc_hd__and2_4
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16411_ _15122_/Y _16406_/X _16410_/X _16406_/X VGND VGND VPWR VPWR _24584_/D sky130_fd_sc_hd__a2bb2o_4
X_13623_ _13623_/A VGND VGND VPWR VPWR _13623_/Y sky130_fd_sc_hd__inv_2
X_17391_ _23973_/Q _20621_/A VGND VGND VPWR VPWR _20625_/A sky130_fd_sc_hd__or2_4
XANTENNA__25094__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_231_0_HCLK clkbuf_8_230_0_HCLK/A VGND VGND VPWR VPWR _24832_/CLK sky130_fd_sc_hd__clkbuf_1
X_19130_ _19130_/A VGND VGND VPWR VPWR _19130_/X sky130_fd_sc_hd__buf_2
XFILLER_73_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16342_ _22478_/A VGND VGND VPWR VPWR _16342_/Y sky130_fd_sc_hd__inv_2
X_13554_ _13554_/A _13554_/B _13550_/X _13553_/X VGND VGND VPWR VPWR _13554_/X sky130_fd_sc_hd__or4_4
XFILLER_12_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25023__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12505_ _12509_/A _12499_/B _12505_/C VGND VGND VPWR VPWR _25421_/D sky130_fd_sc_hd__and3_4
X_19061_ _19105_/A _18331_/X _18922_/X VGND VGND VPWR VPWR _19062_/A sky130_fd_sc_hd__or3_4
X_16273_ _15658_/A _16276_/B VGND VGND VPWR VPWR _16273_/X sky130_fd_sc_hd__or2_4
X_13485_ _13484_/Y _13482_/X _11847_/X _13482_/X VGND VGND VPWR VPWR _13485_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18182__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18012_ _18184_/A _18012_/B _18012_/C VGND VGND VPWR VPWR _18017_/B sky130_fd_sc_hd__and3_4
X_15224_ _15219_/A _15228_/B VGND VGND VPWR VPWR _15225_/C sky130_fd_sc_hd__nand2_4
XFILLER_12_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12436_ _12285_/C _12433_/X VGND VGND VPWR VPWR _12436_/X sky130_fd_sc_hd__or2_4
X_15155_ _15155_/A VGND VGND VPWR VPWR _15155_/Y sky130_fd_sc_hd__inv_2
X_12367_ _12306_/Y _24833_/Q _25342_/Q _12366_/Y VGND VGND VPWR VPWR _12371_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14106_ _14119_/C _14106_/B _14106_/C VGND VGND VPWR VPWR _14107_/C sky130_fd_sc_hd__and3_4
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20661__B2 _17401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12298_ _12377_/A _12296_/Y _13023_/A _24834_/Q VGND VGND VPWR VPWR _12298_/X sky130_fd_sc_hd__a2bb2o_4
X_15086_ _24577_/Q VGND VGND VPWR VPWR _15086_/Y sky130_fd_sc_hd__inv_2
X_19963_ _19963_/A VGND VGND VPWR VPWR _19963_/Y sky130_fd_sc_hd__inv_2
X_14037_ _14012_/A _13999_/X _14010_/C VGND VGND VPWR VPWR _14037_/X sky130_fd_sc_hd__or3_4
X_18914_ _18901_/Y VGND VGND VPWR VPWR _18914_/X sky130_fd_sc_hd__buf_2
XANTENNA__23247__B _22810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19894_ _19894_/A VGND VGND VPWR VPWR _19894_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16617__B1 _16359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18845_ _24539_/Q _18786_/C _24544_/Q _18608_/X VGND VGND VPWR VPWR _18845_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17245__B _17199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24322__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18776_ _18692_/A _18774_/A VGND VGND VPWR VPWR _18776_/X sky130_fd_sc_hd__or2_4
X_15988_ _12231_/Y _15982_/X _15840_/X _15938_/X VGND VGND VPWR VPWR _24736_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12103__B1 _11825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17727_ _24202_/Q VGND VGND VPWR VPWR _17728_/A sky130_fd_sc_hd__buf_2
X_14939_ _14939_/A _14939_/B _14939_/C _14938_/X VGND VGND VPWR VPWR _14939_/X sky130_fd_sc_hd__or4_4
XANTENNA__23958__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_41_0_HCLK clkbuf_6_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_83_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17658_ _17652_/X _17656_/X _17658_/C VGND VGND VPWR VPWR _17658_/X sky130_fd_sc_hd__and3_4
XFILLER_63_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16609_ _16583_/A VGND VGND VPWR VPWR _16609_/X sky130_fd_sc_hd__buf_2
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17589_ _17624_/A VGND VGND VPWR VPWR _17885_/B sky130_fd_sc_hd__inv_2
X_19328_ _19327_/Y _19325_/X _19191_/X _19325_/X VGND VGND VPWR VPWR _23766_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21141__A2 _21335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22607__A _22574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21511__A _21069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19259_ _21373_/B _19256_/X _16888_/X _19256_/X VGND VGND VPWR VPWR _23790_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18092__A _17995_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21429__B1 _11860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22270_ _22646_/A VGND VGND VPWR VPWR _22270_/X sky130_fd_sc_hd__buf_2
X_21221_ _21209_/Y _21103_/X _21211_/X _21220_/X VGND VGND VPWR VPWR _21272_/C sky130_fd_sc_hd__a211o_4
XANTENNA__11749__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24746__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18845__B2 _18608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16856__B1 _16720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21152_ _15670_/A _21149_/X _21151_/X VGND VGND VPWR VPWR _21152_/X sky130_fd_sc_hd__and3_4
X_20103_ _20103_/A VGND VGND VPWR VPWR _22364_/B sky130_fd_sc_hd__inv_2
XANTENNA__12566__A1_N _12565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21083_ _21024_/A VGND VGND VPWR VPWR _22962_/A sky130_fd_sc_hd__buf_2
XFILLER_28_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16340__A HWDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20034_ _21789_/B _20029_/X _19988_/X _20029_/X VGND VGND VPWR VPWR _20034_/X sky130_fd_sc_hd__a2bb2o_4
X_24911_ _24025_/CLK _15558_/X HRESETn VGND VGND VPWR VPWR _23318_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12893__A1 _12841_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_123_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_247_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24842_ _24842_/CLK _15772_/X HRESETn VGND VGND VPWR VPWR _24842_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24773_ _24813_/CLK _15909_/X HRESETn VGND VGND VPWR VPWR _21414_/A sky130_fd_sc_hd__dfrtp_4
X_21985_ _17893_/A _21985_/B VGND VGND VPWR VPWR _21985_/X sky130_fd_sc_hd__and2_4
XANTENNA__13842__B1 _13797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18267__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24107__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25534__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724_ _23722_/CLK _23724_/D VGND VGND VPWR VPWR _23724_/Q sky130_fd_sc_hd__dfxtp_4
X_20936_ _16653_/Y _20814_/X _20909_/A _20935_/Y VGND VGND VPWR VPWR _20936_/X sky130_fd_sc_hd__o22a_4
XPHY_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _24040_/Q VGND VGND VPWR VPWR _20867_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23655_ _24197_/CLK _19654_/X VGND VGND VPWR VPWR _23655_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22606_ _22606_/A VGND VGND VPWR VPWR _22607_/D sky130_fd_sc_hd__inv_2
X_20798_ _20797_/X VGND VGND VPWR VPWR _24024_/D sky130_fd_sc_hd__inv_2
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23586_ _23562_/CLK _19853_/X VGND VGND VPWR VPWR _19851_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25325_ _25351_/CLK _13110_/X HRESETn VGND VGND VPWR VPWR _25325_/Q sky130_fd_sc_hd__dfrtp_4
X_22537_ _22511_/B _22533_/X _22413_/X _22536_/X VGND VGND VPWR VPWR _22537_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_8_61_0_HCLK clkbuf_8_61_0_HCLK/A VGND VGND VPWR VPWR _24712_/CLK sky130_fd_sc_hd__clkbuf_1
X_13270_ _13270_/A _18951_/A VGND VGND VPWR VPWR _13270_/X sky130_fd_sc_hd__or2_4
XANTENNA__20891__B2 _20886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25256_ _24720_/CLK _25256_/D HRESETn VGND VGND VPWR VPWR _25256_/Q sky130_fd_sc_hd__dfrtp_4
X_22468_ _21863_/X _22465_/X _22466_/X _24816_/Q _22467_/X VGND VGND VPWR VPWR _22468_/X
+ sky130_fd_sc_hd__a32o_4
X_12221_ _22465_/A VGND VGND VPWR VPWR _12221_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24487__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24207_ _24214_/CLK _18273_/X HRESETn VGND VGND VPWR VPWR _13695_/A sky130_fd_sc_hd__dfrtp_4
X_21419_ _21418_/X VGND VGND VPWR VPWR _22540_/A sky130_fd_sc_hd__buf_2
X_22399_ _21493_/X _18272_/A _22392_/X _22397_/X _22398_/X VGND VGND VPWR VPWR _22399_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24036__CLK _24581_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21435__A3 _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18836__B2 _18792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25187_ _24942_/CLK _14227_/X HRESETn VGND VGND VPWR VPWR _25187_/Q sky130_fd_sc_hd__dfstp_4
X_12152_ _12152_/A VGND VGND VPWR VPWR _12152_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24416__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24138_ _24136_/CLK _24138_/D HRESETn VGND VGND VPWR VPWR _18603_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_2_2_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12083_ _12083_/A VGND VGND VPWR VPWR _12083_/Y sky130_fd_sc_hd__inv_2
X_16960_ _16960_/A VGND VGND VPWR VPWR _16960_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24069_ _24069_/CLK _20521_/X HRESETn VGND VGND VPWR VPWR _24069_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15911_ _24771_/Q _13590_/A VGND VGND VPWR VPWR _15911_/Y sky130_fd_sc_hd__nor2_4
XFILLER_133_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16891_ _16083_/Y _23314_/A _16083_/Y _23314_/A VGND VGND VPWR VPWR _16895_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17065__B _17260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18630_ _18630_/A VGND VGND VPWR VPWR _18683_/A sky130_fd_sc_hd__inv_2
X_15842_ _15824_/X _15835_/X _15774_/X _24807_/Q _15793_/A VGND VGND VPWR VPWR _24807_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_77_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18561_ _18427_/Y _18580_/A VGND VGND VPWR VPWR _18562_/B sky130_fd_sc_hd__or2_4
XFILLER_76_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15773_ HWDATA[0] VGND VGND VPWR VPWR _15845_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12985_ _25350_/Q VGND VGND VPWR VPWR _13012_/A sky130_fd_sc_hd__inv_2
XFILLER_18_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20500__A _20500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18177__A _18177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25275__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17512_ _17512_/A VGND VGND VPWR VPWR _17512_/Y sky130_fd_sc_hd__inv_2
X_14724_ _14703_/A _14675_/X _14720_/Y _21643_/A _14723_/Y VGND VGND VPWR VPWR _25056_/D
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_5_28_0_HCLK clkbuf_4_14_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_11936_ _11933_/Y _11926_/X _11934_/X _11935_/X VGND VGND VPWR VPWR _25495_/D sky130_fd_sc_hd__a2bb2o_4
X_18492_ _18491_/X VGND VGND VPWR VPWR _18493_/B sky130_fd_sc_hd__inv_2
XANTENNA__25204__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17443_ _17442_/X VGND VGND VPWR VPWR _17443_/X sky130_fd_sc_hd__buf_2
XFILLER_60_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14655_ _14641_/B _14638_/X _14653_/X VGND VGND VPWR VPWR _14655_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15586__B1 _11778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11867_ _11867_/A VGND VGND VPWR VPWR _11867_/X sky130_fd_sc_hd__buf_2
XFILLER_14_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13606_ _13605_/X VGND VGND VPWR VPWR _13606_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12350__A2_N _24821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17374_ _17348_/A _17348_/B _17289_/A _17372_/B VGND VGND VPWR VPWR _17374_/X sky130_fd_sc_hd__a211o_4
X_14586_ _14586_/A VGND VGND VPWR VPWR _14586_/X sky130_fd_sc_hd__buf_2
XANTENNA__17327__A1 _17253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11798_ _25522_/Q VGND VGND VPWR VPWR _11798_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21123__A2 _14220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19113_ _19111_/Y _19107_/X _18997_/X _19112_/X VGND VGND VPWR VPWR _19113_/X sky130_fd_sc_hd__a2bb2o_4
X_16325_ HWDATA[16] VGND VGND VPWR VPWR _16325_/X sky130_fd_sc_hd__buf_2
X_13537_ _13536_/Y _13534_/Y _13472_/X _13534_/Y VGND VGND VPWR VPWR _13537_/X sky130_fd_sc_hd__a2bb2o_4
X_19044_ _19044_/A VGND VGND VPWR VPWR _19044_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16256_ _22089_/A VGND VGND VPWR VPWR _16256_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24064__D _24064_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13468_ _13467_/X VGND VGND VPWR VPWR _13468_/X sky130_fd_sc_hd__buf_2
XFILLER_51_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12365__A2_N _24811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15207_ _15207_/A VGND VGND VPWR VPWR _15207_/Y sky130_fd_sc_hd__inv_2
X_12419_ _12277_/A _12419_/B VGND VGND VPWR VPWR _12420_/C sky130_fd_sc_hd__or2_4
X_16187_ _16187_/A VGND VGND VPWR VPWR _16187_/X sky130_fd_sc_hd__buf_2
X_13399_ _13200_/X _13383_/X _13398_/X _25316_/Q _11964_/X VGND VGND VPWR VPWR _13399_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16838__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15138_ _15369_/A _15122_/A _24984_/Q _15089_/Y VGND VGND VPWR VPWR _15138_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13784__A _16725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17256__A _17247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15069_ _15209_/C _15068_/X VGND VGND VPWR VPWR _15069_/X sky130_fd_sc_hd__or2_4
X_19946_ _19945_/Y _19943_/X _19632_/X _19943_/X VGND VGND VPWR VPWR _19946_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19877_ _23576_/Q VGND VGND VPWR VPWR _21788_/B sky130_fd_sc_hd__inv_2
XFILLER_110_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18828_ _18828_/A _18825_/X _18826_/X _18827_/X VGND VGND VPWR VPWR _18828_/X sky130_fd_sc_hd__or4_4
XFILLER_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13008__B _13008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18759_ _18759_/A _18759_/B _18758_/Y VGND VGND VPWR VPWR _24131_/D sky130_fd_sc_hd__and3_4
XFILLER_23_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13824__B1 _11804_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18087__A _18087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15504__A _15490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21770_ _21623_/A _20054_/Y VGND VGND VPWR VPWR _21770_/X sky130_fd_sc_hd__or2_4
XANTENNA__21225__B _21225_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20721_ _20770_/A VGND VGND VPWR VPWR _20721_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20652_ _14231_/Y _20604_/Y _20619_/A _20651_/X VGND VGND VPWR VPWR _20652_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17535__A1_N _11790_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24998__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23440_ _23441_/CLK _23440_/D VGND VGND VPWR VPWR _13341_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17318__A1 _17254_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12285__D _12433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24927__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23371_ _23904_/CLK _23371_/D VGND VGND VPWR VPWR _23371_/Q sky130_fd_sc_hd__dfxtp_4
X_20583_ _18880_/X VGND VGND VPWR VPWR _20583_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_48_0_HCLK clkbuf_6_24_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_48_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_25110_ _23959_/CLK _25110_/D HRESETn VGND VGND VPWR VPWR _25110_/Q sky130_fd_sc_hd__dfrtp_4
X_22322_ _22321_/X VGND VGND VPWR VPWR _22322_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13678__B _13678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_5_19_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22253_ _21478_/A _22253_/B VGND VGND VPWR VPWR _22254_/C sky130_fd_sc_hd__or2_4
XANTENNA__24580__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25041_ _25043_/CLK _25041_/D HRESETn VGND VGND VPWR VPWR _14803_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_3_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21204_ _24310_/Q _13782_/A VGND VGND VPWR VPWR _21204_/X sky130_fd_sc_hd__and2_4
XFILLER_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22184_ _21859_/B _22183_/X _21284_/A VGND VGND VPWR VPWR _22184_/X sky130_fd_sc_hd__and3_4
XANTENNA__22072__A _21618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21135_ _21014_/A _21135_/B VGND VGND VPWR VPWR _21135_/Y sky130_fd_sc_hd__nor2_4
XFILLER_105_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21066_ _21066_/A VGND VGND VPWR VPWR _21067_/A sky130_fd_sc_hd__buf_2
XFILLER_24_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20389__B1 _15766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20017_ _20016_/Y _20014_/X _19995_/X _20014_/X VGND VGND VPWR VPWR _23526_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21416__A _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24825_ _24852_/CLK _24825_/D HRESETn VGND VGND VPWR VPWR _24825_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17006__B1 _24731_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12770_ _25363_/Q _24780_/Q _12944_/B _12769_/Y VGND VGND VPWR VPWR _12777_/B sky130_fd_sc_hd__o22a_4
XFILLER_73_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24756_ _24759_/CLK _15956_/X HRESETn VGND VGND VPWR VPWR _22964_/A sky130_fd_sc_hd__dfrtp_4
X_21968_ _21968_/A _20318_/X VGND VGND VPWR VPWR _21968_/X sky130_fd_sc_hd__or2_4
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21353__A2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18754__B1 _18707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _16079_/A VGND VGND VPWR VPWR _11739_/A sky130_fd_sc_hd__inv_2
XANTENNA__14675__D _13593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _23598_/CLK _23707_/D VGND VGND VPWR VPWR _23707_/Q sky130_fd_sc_hd__dfxtp_4
X_20919_ _20918_/Y _20915_/Y _20922_/B VGND VGND VPWR VPWR _20919_/X sky130_fd_sc_hd__o21a_4
XPHY_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24687_ _24689_/CLK _16119_/X HRESETn VGND VGND VPWR VPWR _22902_/A sky130_fd_sc_hd__dfrtp_4
X_21899_ _14689_/A _21899_/B VGND VGND VPWR VPWR _21901_/B sky130_fd_sc_hd__or2_4
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14439_/Y _14437_/X _14414_/X _14437_/X VGND VGND VPWR VPWR _25123_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _21504_/A _11970_/C VGND VGND VPWR VPWR _11652_/X sky130_fd_sc_hd__and2_4
XFILLER_70_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23638_ _24288_/CLK _23638_/D VGND VGND VPWR VPWR _19699_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_70_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14240__B1 _14239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24668__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ _14354_/Y _14370_/X _12088_/A _14330_/X VGND VGND VPWR VPWR _14371_/X sky130_fd_sc_hd__o22a_4
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23569_ _23545_/CLK _19898_/X VGND VGND VPWR VPWR _19897_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_31_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16110_ _24690_/Q VGND VGND VPWR VPWR _16110_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13322_ _13390_/A _13322_/B _13321_/X VGND VGND VPWR VPWR _13333_/B sky130_fd_sc_hd__or3_4
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25308_ _25305_/CLK _13485_/X HRESETn VGND VGND VPWR VPWR _13484_/A sky130_fd_sc_hd__dfrtp_4
X_17090_ _17020_/X VGND VGND VPWR VPWR _17108_/A sky130_fd_sc_hd__buf_2
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16041_ _16039_/Y _16035_/X _11804_/X _16040_/X VGND VGND VPWR VPWR _24717_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13253_ _13395_/A _13253_/B VGND VGND VPWR VPWR _13253_/X sky130_fd_sc_hd__or2_4
X_25239_ _24148_/CLK _13865_/X HRESETn VGND VGND VPWR VPWR _20466_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12204_ _24743_/Q VGND VGND VPWR VPWR _12204_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24250__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_5_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__21813__B1 _21679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13184_ _13188_/A _13182_/X _13183_/X VGND VGND VPWR VPWR _13184_/X sky130_fd_sc_hd__and3_4
XFILLER_124_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19800_ _21229_/B _19793_/X _18919_/X _19793_/A VGND VGND VPWR VPWR _23605_/D sky130_fd_sc_hd__a2bb2o_4
X_12135_ _12113_/A _12134_/A _12113_/Y _12134_/Y VGND VGND VPWR VPWR _12135_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17493__B1 _11706_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17992_ _18181_/A _17992_/B _17992_/C VGND VGND VPWR VPWR _17993_/C sky130_fd_sc_hd__and3_4
XFILLER_97_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16943_ _24267_/Q VGND VGND VPWR VPWR _16943_/Y sky130_fd_sc_hd__inv_2
X_19731_ _19727_/Y _19730_/X _19664_/X _19730_/X VGND VGND VPWR VPWR _23628_/D sky130_fd_sc_hd__a2bb2o_4
X_12066_ _21559_/A VGND VGND VPWR VPWR _12066_/X sky130_fd_sc_hd__buf_2
XFILLER_78_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21041__A1 _24842_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25456__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19291__A _19642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16874_ _20092_/A VGND VGND VPWR VPWR _19790_/A sky130_fd_sc_hd__buf_2
X_19662_ _19661_/X VGND VGND VPWR VPWR _19676_/A sky130_fd_sc_hd__inv_2
XFILLER_64_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15825_ _15824_/X _15819_/X _11818_/A _24818_/Q _15793_/A VGND VGND VPWR VPWR _24818_/D
+ sky130_fd_sc_hd__a32o_4
X_18613_ _24523_/Q _18749_/A _24529_/Q _18696_/A VGND VGND VPWR VPWR _18616_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21326__A _22798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19593_ _19587_/X VGND VGND VPWR VPWR _19593_/X sky130_fd_sc_hd__buf_2
XANTENNA__15953__A1_N _12259_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11852__A _18254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15756_ HWDATA[9] VGND VGND VPWR VPWR _15756_/X sky130_fd_sc_hd__buf_2
X_18544_ _18532_/B VGND VGND VPWR VPWR _18545_/B sky130_fd_sc_hd__inv_2
X_12968_ _12819_/X _12941_/X _12884_/A _12966_/B VGND VGND VPWR VPWR _12969_/A sky130_fd_sc_hd__a211o_4
XFILLER_92_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22541__A1 _24544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14707_ _14707_/A VGND VGND VPWR VPWR _14707_/Y sky130_fd_sc_hd__inv_2
X_11919_ _11902_/B _11910_/X VGND VGND VPWR VPWR _11919_/Y sky130_fd_sc_hd__nor2_4
X_18475_ _18427_/Y _18475_/B _18475_/C _18475_/D VGND VGND VPWR VPWR _18476_/C sky130_fd_sc_hd__or4_4
XFILLER_33_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15687_ _15687_/A _15687_/B _15687_/C VGND VGND VPWR VPWR _15687_/X sky130_fd_sc_hd__or3_4
X_12899_ _12882_/A _12896_/B _12898_/X VGND VGND VPWR VPWR _12900_/A sky130_fd_sc_hd__or3_4
X_17426_ _17423_/Y _17417_/X _17424_/X _17425_/X VGND VGND VPWR VPWR _17426_/X sky130_fd_sc_hd__a2bb2o_4
X_14638_ _14620_/D _13633_/B _13635_/A VGND VGND VPWR VPWR _14638_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21061__A _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17357_ _17357_/A VGND VGND VPWR VPWR _17357_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14569_ _14569_/A VGND VGND VPWR VPWR _14570_/B sky130_fd_sc_hd__inv_2
XANTENNA__19170__B1 _19056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16308_ _23009_/A VGND VGND VPWR VPWR _16308_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24338__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17288_ _17258_/B _17267_/X _17236_/Y VGND VGND VPWR VPWR _17288_/X sky130_fd_sc_hd__o21a_4
XFILLER_101_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19027_ _23872_/Q VGND VGND VPWR VPWR _19027_/Y sky130_fd_sc_hd__inv_2
X_16239_ _16237_/Y _16232_/X _16238_/X _16232_/X VGND VGND VPWR VPWR _16239_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15994__A _22915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15731__B1 _11774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20607__A1 _14868_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14403__A _16359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19929_ _19929_/A VGND VGND VPWR VPWR _19929_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23973__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25197__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22940_ _22940_/A _22394_/X _22812_/C VGND VGND VPWR VPWR _22940_/X sky130_fd_sc_hd__and3_4
XFILLER_56_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22780__B2 _22288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20140__A _20140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22871_ _22869_/X _22870_/X _22440_/C VGND VGND VPWR VPWR _22871_/X sky130_fd_sc_hd__or3_4
X_24610_ _24177_/CLK _24610_/D HRESETn VGND VGND VPWR VPWR _16336_/A sky130_fd_sc_hd__dfrtp_4
X_21822_ _21815_/Y _21821_/X _22035_/A VGND VGND VPWR VPWR _21822_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18848__A1_N _24551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_11_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24541_ _24541_/CLK _24541_/D HRESETn VGND VGND VPWR VPWR _24541_/Q sky130_fd_sc_hd__dfrtp_4
X_21753_ _21608_/A _21753_/B VGND VGND VPWR VPWR _21753_/X sky130_fd_sc_hd__or2_4
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20704_ _22281_/A _20698_/X _20686_/X _20703_/Y VGND VGND VPWR VPWR _20704_/X sky130_fd_sc_hd__o22a_4
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24472_ _24649_/CLK _24472_/D HRESETn VGND VGND VPWR VPWR _24472_/Q sky130_fd_sc_hd__dfrtp_4
X_21684_ _13795_/D _21683_/X _18265_/A _18261_/A VGND VGND VPWR VPWR _21684_/X sky130_fd_sc_hd__o22a_4
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22067__A _14682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21099__A1 _17242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22296__B1 _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24761__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23423_ _24923_/CLK _20288_/X VGND VGND VPWR VPWR _23423_/Q sky130_fd_sc_hd__dfxtp_4
X_20635_ _20638_/B _20635_/B _20651_/C VGND VGND VPWR VPWR _20635_/X sky130_fd_sc_hd__and3_4
XFILLER_123_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15970__B1 _24750_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19161__B1 _19136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24079__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20566_ _20566_/A _20566_/B VGND VGND VPWR VPWR _20567_/B sky130_fd_sc_hd__nand2_4
X_23354_ _23338_/X VGND VGND VPWR VPWR IRQ[0] sky130_fd_sc_hd__buf_2
XFILLER_20_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24008__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22305_ _14381_/A _17415_/A _25096_/Q _22172_/B VGND VGND VPWR VPWR _22309_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25087__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15722__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20497_ _14386_/A _14495_/X _20495_/X _20457_/D _20496_/X VGND VGND VPWR VPWR _20497_/X
+ sky130_fd_sc_hd__a32o_4
X_23285_ _23285_/A _23226_/B VGND VGND VPWR VPWR _23285_/X sky130_fd_sc_hd__and2_4
XANTENNA__22599__A1 _21105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25024_ _25024_/CLK _25024_/D HRESETn VGND VGND VPWR VPWR _15179_/A sky130_fd_sc_hd__dfrtp_4
X_22236_ _22247_/A _22234_/X _22235_/X VGND VGND VPWR VPWR _22236_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_135_0_HCLK clkbuf_7_67_0_HCLK/X VGND VGND VPWR VPWR _23904_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_3_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21271__A1 _21261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_198_0_HCLK clkbuf_7_99_0_HCLK/X VGND VGND VPWR VPWR _24026_/CLK sky130_fd_sc_hd__clkbuf_1
X_22167_ _21826_/A _22166_/X VGND VGND VPWR VPWR _22167_/X sky130_fd_sc_hd__and2_4
X_21118_ _21143_/A VGND VGND VPWR VPWR _21333_/A sky130_fd_sc_hd__inv_2
XFILLER_59_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22098_ _22097_/Y _21336_/A _14416_/Y _21338_/X VGND VGND VPWR VPWR _22098_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22530__A _22574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13940_ _13939_/X VGND VGND VPWR VPWR _13970_/A sky130_fd_sc_hd__inv_2
X_21049_ _22913_/A VGND VGND VPWR VPWR _21049_/X sky130_fd_sc_hd__buf_2
XANTENNA__17624__A _17624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18975__B1 _18955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20945__A1_N _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13871_ _23989_/Q VGND VGND VPWR VPWR _13871_/X sky130_fd_sc_hd__buf_2
X_15610_ _15609_/Y _15605_/X _11818_/X _15605_/X VGND VGND VPWR VPWR _24891_/D sky130_fd_sc_hd__a2bb2o_4
X_12822_ _24792_/Q VGND VGND VPWR VPWR _12822_/Y sky130_fd_sc_hd__inv_2
X_24808_ _24836_/CLK _24808_/D HRESETn VGND VGND VPWR VPWR _24808_/Q sky130_fd_sc_hd__dfrtp_4
X_16590_ _16590_/A VGND VGND VPWR VPWR _16590_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15541_ _15540_/Y _15538_/X HADDR[1] _15538_/X VGND VGND VPWR VPWR _15541_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23361__A _21004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24849__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12753_ _12753_/A VGND VGND VPWR VPWR _12753_/X sky130_fd_sc_hd__buf_2
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24739_ _24766_/CLK _15984_/X HRESETn VGND VGND VPWR VPWR _24739_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14983__A _14976_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11704_/A VGND VGND VPWR VPWR _11967_/C sky130_fd_sc_hd__inv_2
X_18260_ _13791_/X VGND VGND VPWR VPWR _18261_/A sky130_fd_sc_hd__buf_2
XFILLER_30_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _15470_/Y _15468_/X _15471_/X _15468_/X VGND VGND VPWR VPWR _15472_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12686_/A _12684_/B _12683_/Y VGND VGND VPWR VPWR _25405_/D sky130_fd_sc_hd__and3_4
XANTENNA__14213__B1 _13515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23079__A2 _22824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17204_/X _17211_/B _17211_/C _17211_/D VGND VGND VPWR VPWR _17230_/A sky130_fd_sc_hd__or4_4
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _25128_/Q VGND VGND VPWR VPWR _14423_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13599__A _13598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18191_ _18191_/A _18189_/X _18190_/X VGND VGND VPWR VPWR _18192_/C sky130_fd_sc_hd__and3_4
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15961__B1 _15959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17142_ _17038_/B _17132_/X VGND VGND VPWR VPWR _17143_/C sky130_fd_sc_hd__nand2_4
XANTENNA__24431__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14354_ _14330_/X VGND VGND VPWR VPWR _14354_/Y sky130_fd_sc_hd__inv_2
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22705__A _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13305_ _13301_/X _13303_/X _13305_/C VGND VGND VPWR VPWR _13305_/X sky130_fd_sc_hd__and3_4
XFILLER_13_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_31_0_HCLK clkbuf_7_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17073_ _17064_/A _17073_/B _17072_/X VGND VGND VPWR VPWR _17073_/X sky130_fd_sc_hd__and3_4
X_14285_ _23428_/Q _14280_/X _14283_/X _25171_/Q _14284_/Y VGND VGND VPWR VPWR _25171_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_7_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18190__A _18046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_94_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_94_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16024_ _24723_/Q VGND VGND VPWR VPWR _16024_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13236_ _13227_/A VGND VGND VPWR VPWR _13317_/A sky130_fd_sc_hd__buf_2
XFILLER_108_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11847__A _16355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13167_ _13188_/A _13164_/X _13166_/X VGND VGND VPWR VPWR _13167_/X sky130_fd_sc_hd__and3_4
X_12118_ _25458_/Q VGND VGND VPWR VPWR _12118_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13098_ _12377_/Y _13082_/X VGND VGND VPWR VPWR _13100_/B sky130_fd_sc_hd__nand2_4
X_17975_ _17975_/A VGND VGND VPWR VPWR _17990_/A sky130_fd_sc_hd__buf_2
XANTENNA__25290__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_0_0_HCLK clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19714_ _23633_/Q VGND VGND VPWR VPWR _19714_/Y sky130_fd_sc_hd__inv_2
X_12049_ _12049_/A VGND VGND VPWR VPWR _12050_/A sky130_fd_sc_hd__inv_2
X_16926_ _16926_/A VGND VGND VPWR VPWR _16927_/A sky130_fd_sc_hd__inv_2
XFILLER_84_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14976__A2_N _16850_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18966__B1 _17443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19645_ _18996_/X VGND VGND VPWR VPWR _19645_/X sky130_fd_sc_hd__buf_2
X_16857_ _20079_/A VGND VGND VPWR VPWR _19777_/A sky130_fd_sc_hd__buf_2
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15808_ _12368_/Y _15802_/X _11774_/X _15802_/X VGND VGND VPWR VPWR _15808_/X sky130_fd_sc_hd__a2bb2o_4
X_16788_ _16785_/Y _16783_/X _16787_/X _16783_/X VGND VGND VPWR VPWR _16788_/X sky130_fd_sc_hd__a2bb2o_4
X_19576_ _19576_/A VGND VGND VPWR VPWR _19576_/Y sky130_fd_sc_hd__inv_2
X_15739_ HWDATA[16] VGND VGND VPWR VPWR _15739_/X sky130_fd_sc_hd__buf_2
X_18527_ _18400_/Y _18525_/A VGND VGND VPWR VPWR _18527_/X sky130_fd_sc_hd__or2_4
XANTENNA__21868__A3 _22644_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24519__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18458_ _24168_/Q VGND VGND VPWR VPWR _18458_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14204__B1 _13837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17409_ _17387_/X _17401_/X _20990_/B _24323_/Q _17404_/X VGND VGND VPWR VPWR _24323_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_5_0_HCLK_A clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18389_ _24631_/Q VGND VGND VPWR VPWR _18389_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22817__A2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15830__A1_N _12318_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20420_ _25138_/Q _20420_/B VGND VGND VPWR VPWR _20421_/A sky130_fd_sc_hd__or2_4
XANTENNA__13302__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24172__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24101__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20351_ _20351_/A VGND VGND VPWR VPWR _21654_/B sky130_fd_sc_hd__inv_2
XANTENNA__16613__A _24506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23070_ _24526_/Q _22393_/X _15668_/A _23069_/X VGND VGND VPWR VPWR _23071_/C sky130_fd_sc_hd__a211o_4
X_20282_ _23425_/Q VGND VGND VPWR VPWR _22006_/B sky130_fd_sc_hd__inv_2
XFILLER_127_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22021_ _22024_/A _19520_/Y VGND VGND VPWR VPWR _22021_/X sky130_fd_sc_hd__or2_4
XANTENNA__25378__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11757__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_208_0_HCLK clkbuf_7_104_0_HCLK/X VGND VGND VPWR VPWR _24496_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25307__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23972_ _24943_/CLK _23972_/D HRESETn VGND VGND VPWR VPWR _20620_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_111_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22923_ _22923_/A VGND VGND VPWR VPWR _22923_/X sky130_fd_sc_hd__buf_2
XANTENNA__20764__B1 _20706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22854_ _22466_/A VGND VGND VPWR VPWR _22854_/X sky130_fd_sc_hd__buf_2
XANTENNA__14443__B1 _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21805_ _21671_/A _21803_/X _21804_/X VGND VGND VPWR VPWR _21805_/X sky130_fd_sc_hd__and3_4
XANTENNA__12100__B _13496_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22785_ _16680_/Y _22872_/B VGND VGND VPWR VPWR _22785_/X sky130_fd_sc_hd__and2_4
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19382__B1 _19291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24524_ _24557_/CLK _16568_/X HRESETn VGND VGND VPWR VPWR _24524_/Q sky130_fd_sc_hd__dfrtp_4
X_21736_ _22441_/A _21733_/X _22444_/A _21735_/X VGND VGND VPWR VPWR _21737_/B sky130_fd_sc_hd__o22a_4
XANTENNA__16196__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22269__B1 _12296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24455_ _25024_/CLK _16748_/X HRESETn VGND VGND VPWR VPWR _24455_/Q sky130_fd_sc_hd__dfrtp_4
X_21667_ _21191_/A VGND VGND VPWR VPWR _21668_/A sky130_fd_sc_hd__buf_2
XANTENNA__15943__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19134__B1 _19133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20819__A1 _16719_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23406_ _24208_/CLK _23406_/D VGND VGND VPWR VPWR _20331_/A sky130_fd_sc_hd__dfxtp_4
X_20618_ _14807_/A VGND VGND VPWR VPWR _20619_/A sky130_fd_sc_hd__buf_2
XANTENNA__20819__B2 _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24386_ _24391_/CLK _17076_/Y HRESETn VGND VGND VPWR VPWR _17026_/A sky130_fd_sc_hd__dfrtp_4
X_21598_ _21630_/A _21598_/B VGND VGND VPWR VPWR _21599_/C sky130_fd_sc_hd__or2_4
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22525__A _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_18_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_18_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23337_ _13799_/A _21964_/X _23335_/Y _23336_/Y VGND VGND VPWR VPWR _23337_/X sky130_fd_sc_hd__a211o_4
X_20549_ _18873_/B _20548_/Y _20558_/C VGND VGND VPWR VPWR _20549_/X sky130_fd_sc_hd__and3_4
XANTENNA__16523__A _24540_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14070_ _14070_/A _14070_/B VGND VGND VPWR VPWR _14071_/B sky130_fd_sc_hd__or2_4
X_23268_ _23245_/X _23249_/X _23268_/C _23267_/X VGND VGND VPWR VPWR HRDATA[29] sky130_fd_sc_hd__or4_4
X_13021_ _13023_/B VGND VGND VPWR VPWR _13026_/B sky130_fd_sc_hd__inv_2
X_25007_ _25010_/CLK _15245_/Y HRESETn VGND VGND VPWR VPWR _14947_/A sky130_fd_sc_hd__dfrtp_4
X_22219_ _14716_/A _22211_/X _22218_/X VGND VGND VPWR VPWR _22219_/X sky130_fd_sc_hd__and3_4
X_23199_ _23128_/A _23199_/B VGND VGND VPWR VPWR _23199_/Y sky130_fd_sc_hd__nor2_4
XFILLER_121_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25048__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23356__A _23343_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14972_ _25015_/Q VGND VGND VPWR VPWR _15212_/A sky130_fd_sc_hd__inv_2
X_17760_ _17751_/X _17760_/B VGND VGND VPWR VPWR _17792_/B sky130_fd_sc_hd__or2_4
XFILLER_0_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18948__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22744__B2 _22743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13923_ _13919_/X _13920_/X _13889_/C _24954_/Q VGND VGND VPWR VPWR _13930_/B sky130_fd_sc_hd__a211o_4
X_16711_ _16711_/A VGND VGND VPWR VPWR _16711_/Y sky130_fd_sc_hd__inv_2
X_17691_ _17662_/A _17689_/X VGND VGND VPWR VPWR _17691_/X sky130_fd_sc_hd__or2_4
XANTENNA__12498__A _12280_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16642_ _24496_/Q VGND VGND VPWR VPWR _23285_/A sky130_fd_sc_hd__inv_2
X_19430_ _18034_/B VGND VGND VPWR VPWR _19430_/Y sky130_fd_sc_hd__inv_2
X_13854_ _13853_/A _13851_/X _13852_/X _13853_/Y VGND VGND VPWR VPWR _25241_/D sky130_fd_sc_hd__a211o_4
XFILLER_63_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12805_ _25368_/Q VGND VGND VPWR VPWR _12806_/A sky130_fd_sc_hd__inv_2
XANTENNA__20899__A1_N _20882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24683__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16573_ _16572_/Y _16570_/X _16403_/X _16570_/X VGND VGND VPWR VPWR _24522_/D sky130_fd_sc_hd__a2bb2o_4
X_19361_ _19355_/Y VGND VGND VPWR VPWR _19361_/X sky130_fd_sc_hd__buf_2
XFILLER_16_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13785_ _13770_/X _13784_/X _13472_/X _13784_/X VGND VGND VPWR VPWR _13785_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19373__B1 _19349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15524_ _15535_/A VGND VGND VPWR VPWR _15524_/X sky130_fd_sc_hd__buf_2
X_18312_ _24202_/Q VGND VGND VPWR VPWR _21196_/A sky130_fd_sc_hd__inv_2
XANTENNA__24612__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12736_ _25389_/Q _12736_/B VGND VGND VPWR VPWR _12736_/X sky130_fd_sc_hd__or2_4
X_19292_ _19290_/Y _19288_/X _19291_/X _19288_/X VGND VGND VPWR VPWR _23779_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18243_ _11671_/Y _18233_/X _15752_/X _18242_/X VGND VGND VPWR VPWR _24224_/D sky130_fd_sc_hd__a2bb2o_4
X_15455_ _13895_/X _15449_/X _15446_/X _24950_/Q _15452_/X VGND VGND VPWR VPWR _15455_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_54_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12667_ _12611_/B _12666_/X VGND VGND VPWR VPWR _12670_/B sky130_fd_sc_hd__or2_4
XANTENNA__15934__B1 _24766_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ _14406_/A _18895_/A VGND VGND VPWR VPWR _14407_/A sky130_fd_sc_hd__or2_4
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18174_ _17973_/X _19461_/A VGND VGND VPWR VPWR _18174_/X sky130_fd_sc_hd__or2_4
XFILLER_50_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15386_ _15385_/X VGND VGND VPWR VPWR _15386_/Y sky130_fd_sc_hd__inv_2
X_12598_ _12598_/A _12593_/X _12598_/C _12598_/D VGND VGND VPWR VPWR _12598_/X sky130_fd_sc_hd__or4_4
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17125_ _17120_/A _17119_/X _17121_/Y _17056_/X VGND VGND VPWR VPWR _17126_/A sky130_fd_sc_hd__a211o_4
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14337_ _25151_/Q VGND VGND VPWR VPWR _14337_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22154__B _22298_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17056_ _17384_/B VGND VGND VPWR VPWR _17056_/X sky130_fd_sc_hd__buf_2
XANTENNA__15029__A2_N _15027_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14268_ _14268_/A VGND VGND VPWR VPWR _14268_/Y sky130_fd_sc_hd__inv_2
X_16007_ _24730_/Q VGND VGND VPWR VPWR _16007_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25471__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13219_ _13225_/A VGND VGND VPWR VPWR _13269_/A sky130_fd_sc_hd__buf_2
X_14199_ _14210_/B _14196_/X _14200_/A VGND VGND VPWR VPWR _14199_/X sky130_fd_sc_hd__a21o_4
XFILLER_112_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25400__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16111__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_181_0_HCLK clkbuf_7_90_0_HCLK/X VGND VGND VPWR VPWR _24692_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_38_0_HCLK clkbuf_8_39_0_HCLK/A VGND VGND VPWR VPWR _25044_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17958_ _17954_/X _17957_/X _18006_/A VGND VGND VPWR VPWR _17958_/X sky130_fd_sc_hd__o21a_4
XFILLER_100_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16909_ _24269_/Q VGND VGND VPWR VPWR _16909_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20746__B1 _20745_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17889_ _17891_/A VGND VGND VPWR VPWR _17889_/X sky130_fd_sc_hd__buf_2
XFILLER_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24938__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19628_ _19628_/A VGND VGND VPWR VPWR _19628_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19559_ _23684_/Q VGND VGND VPWR VPWR _22342_/B sky130_fd_sc_hd__inv_2
XFILLER_20_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16608__A _16608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24353__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22570_ _22530_/X _22538_/Y _22543_/X _22570_/D VGND VGND VPWR VPWR HRDATA[10] sky130_fd_sc_hd__or4_4
XFILLER_55_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21521_ _21512_/X _21519_/X _21514_/X _12552_/A _21520_/X VGND VGND VPWR VPWR _21521_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_33_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18823__A pwm_S7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24240_ _23805_/CLK _24240_/D HRESETn VGND VGND VPWR VPWR _17911_/A sky130_fd_sc_hd__dfrtp_4
X_21452_ _21452_/A _21449_/X _21451_/X VGND VGND VPWR VPWR _21452_/X sky130_fd_sc_hd__and3_4
XFILLER_33_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20403_ _20402_/Y _20400_/X _19755_/X _20400_/X VGND VGND VPWR VPWR _23377_/D sky130_fd_sc_hd__a2bb2o_4
X_21383_ _21398_/A _21381_/X _21383_/C VGND VGND VPWR VPWR _21383_/X sky130_fd_sc_hd__and3_4
X_24171_ _24171_/CLK _24171_/D HRESETn VGND VGND VPWR VPWR _24171_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23122_ _15574_/Y _23052_/B VGND VGND VPWR VPWR _23122_/X sky130_fd_sc_hd__and2_4
X_20334_ _21985_/B _20327_/X _18267_/X _20326_/Y VGND VGND VPWR VPWR _23405_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20265_ _20265_/A VGND VGND VPWR VPWR _21626_/B sky130_fd_sc_hd__inv_2
XANTENNA__22423__B1 _16054_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23053_ _22783_/X _23051_/X _22786_/X _23052_/X VGND VGND VPWR VPWR _23053_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21777__A2 _21776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25141__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22004_ _22016_/A _22004_/B VGND VGND VPWR VPWR _22007_/B sky130_fd_sc_hd__or2_4
XANTENNA__16102__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20196_ _20203_/A VGND VGND VPWR VPWR _20196_/X sky130_fd_sc_hd__buf_2
XFILLER_89_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20985__B1 _20490_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23955_ _24318_/CLK _23955_/D HRESETn VGND VGND VPWR VPWR _23955_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_9_0_HCLK clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__17602__B1 _17601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22906_ _22186_/A VGND VGND VPWR VPWR _22906_/X sky130_fd_sc_hd__buf_2
X_23886_ _23887_/CLK _23886_/D VGND VGND VPWR VPWR _18982_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21424__A _21071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22837_ _24418_/Q _22833_/X _22834_/X _22836_/X VGND VGND VPWR VPWR _22838_/C sky130_fd_sc_hd__a211o_4
XFILLER_32_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24094__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ _13570_/A VGND VGND VPWR VPWR _13570_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22768_ _22897_/A _22768_/B VGND VGND VPWR VPWR _22778_/C sky130_fd_sc_hd__and2_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _12520_/Y VGND VGND VPWR VPWR _12679_/A sky130_fd_sc_hd__buf_2
XFILLER_72_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24023__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24507_ _24541_/CLK _24507_/D HRESETn VGND VGND VPWR VPWR _16611_/A sky130_fd_sc_hd__dfrtp_4
X_21719_ _14216_/Y _14194_/A _14233_/Y _21338_/X VGND VGND VPWR VPWR _21720_/A sky130_fd_sc_hd__o22a_4
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25487_ _23384_/CLK _11971_/Y HRESETn VGND VGND VPWR VPWR _11967_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__18664__A1_N _24530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22699_ _16503_/A _22695_/B _21859_/C VGND VGND VPWR VPWR _22699_/X sky130_fd_sc_hd__and3_4
XFILLER_40_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A VGND VGND VPWR VPWR _15240_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12452_ _12238_/X _12430_/X VGND VGND VPWR VPWR _12455_/B sky130_fd_sc_hd__or2_4
X_24438_ _24407_/CLK _24438_/D HRESETn VGND VGND VPWR VPWR _14991_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15171_ _14986_/A _15171_/B VGND VGND VPWR VPWR _15171_/X sky130_fd_sc_hd__and2_4
X_12383_ _12382_/X VGND VGND VPWR VPWR _13008_/B sky130_fd_sc_hd__buf_2
XFILLER_123_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24369_ _24364_/CLK _24369_/D HRESETn VGND VGND VPWR VPWR _16983_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25229__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14122_ _23950_/Q VGND VGND VPWR VPWR _14181_/B sky130_fd_sc_hd__buf_2
XFILLER_126_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16341__B1 _16340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23206__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14053_ _14012_/A _14047_/Y _14010_/C VGND VGND VPWR VPWR _14053_/X sky130_fd_sc_hd__or3_4
X_18930_ _18937_/A VGND VGND VPWR VPWR _18930_/X sky130_fd_sc_hd__buf_2
XFILLER_137_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13004_ _25353_/Q _13004_/B VGND VGND VPWR VPWR _13004_/X sky130_fd_sc_hd__or2_4
XFILLER_97_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22702__B _21220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18861_ _16457_/Y _18599_/X _16457_/Y _18599_/X VGND VGND VPWR VPWR _18861_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18602__A1_N _16608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_254_0_HCLK clkbuf_8_255_0_HCLK/A VGND VGND VPWR VPWR _25411_/CLK sky130_fd_sc_hd__clkbuf_1
X_17812_ _17814_/B VGND VGND VPWR VPWR _17813_/B sky130_fd_sc_hd__inv_2
XFILLER_121_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18792_ _18792_/A _18792_/B _18792_/C VGND VGND VPWR VPWR _18792_/X sky130_fd_sc_hd__or3_4
X_14955_ _25018_/Q VGND VGND VPWR VPWR _14955_/Y sky130_fd_sc_hd__inv_2
X_17743_ _17743_/A _16909_/Y VGND VGND VPWR VPWR _17761_/C sky130_fd_sc_hd__or2_4
XANTENNA__15316__B _15165_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24864__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19594__B1 _19407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13906_ _13909_/C _24950_/Q _13899_/X _13905_/B VGND VGND VPWR VPWR _13906_/X sky130_fd_sc_hd__or4_4
X_14886_ _14885_/Y VGND VGND VPWR VPWR _14886_/X sky130_fd_sc_hd__buf_2
X_17674_ _17517_/Y _17674_/B VGND VGND VPWR VPWR _17675_/C sky130_fd_sc_hd__nand2_4
XFILLER_36_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19413_ _19412_/Y _19408_/X _19389_/X _19408_/X VGND VGND VPWR VPWR _19413_/X sky130_fd_sc_hd__a2bb2o_4
X_13837_ _11838_/A VGND VGND VPWR VPWR _13837_/X sky130_fd_sc_hd__buf_2
X_16625_ _16624_/X VGND VGND VPWR VPWR _16625_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22149__B _22149_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11860__A _11860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16556_ _16555_/Y _16551_/X _16386_/X _16551_/X VGND VGND VPWR VPWR _16556_/X sky130_fd_sc_hd__a2bb2o_4
X_19344_ _19343_/Y _19339_/X _19232_/X _19339_/X VGND VGND VPWR VPWR _19344_/X sky130_fd_sc_hd__a2bb2o_4
X_13768_ _13748_/A _14703_/A _20043_/D VGND VGND VPWR VPWR _25264_/D sky130_fd_sc_hd__o21a_4
X_12719_ _12698_/A _12707_/B _12719_/C VGND VGND VPWR VPWR _25395_/D sky130_fd_sc_hd__and3_4
X_15507_ _15506_/Y _15504_/X HADDR[16] _15504_/X VGND VGND VPWR VPWR _15507_/X sky130_fd_sc_hd__a2bb2o_4
X_16487_ _16485_/Y _16486_/X _16401_/X _16486_/X VGND VGND VPWR VPWR _16487_/X sky130_fd_sc_hd__a2bb2o_4
X_19275_ _23784_/Q VGND VGND VPWR VPWR _21752_/B sky130_fd_sc_hd__inv_2
XANTENNA__15907__B1 _24775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13699_ _13702_/A _13702_/B VGND VGND VPWR VPWR _13699_/X sky130_fd_sc_hd__or2_4
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15438_ _15434_/X VGND VGND VPWR VPWR _15438_/X sky130_fd_sc_hd__buf_2
X_18226_ _15694_/X _18210_/X _18225_/X _24230_/Q _18019_/A VGND VGND VPWR VPWR _18226_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__16580__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12197__B2 _24735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15369_ _15369_/A _15369_/B VGND VGND VPWR VPWR _15370_/C sky130_fd_sc_hd__nand2_4
X_18157_ _18054_/X _19187_/A VGND VGND VPWR VPWR _18159_/B sky130_fd_sc_hd__or2_4
XANTENNA__17259__A _17178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18321__A1 _24198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17108_ _17108_/A _17108_/B _17107_/Y VGND VGND VPWR VPWR _24378_/D sky130_fd_sc_hd__and3_4
XFILLER_89_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18088_ _18088_/A VGND VGND VPWR VPWR _18186_/A sky130_fd_sc_hd__buf_2
XFILLER_132_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17039_ _17039_/A VGND VGND VPWR VPWR _17156_/A sky130_fd_sc_hd__inv_2
XFILLER_116_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20050_ _20057_/A VGND VGND VPWR VPWR _20050_/X sky130_fd_sc_hd__buf_2
XFILLER_113_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14411__A _16057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15989__A3 _15927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20719__B1 _20706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18388__A1 _24103_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15536__A2_N _15535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17722__A _17722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24534__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23740_ _23828_/CLK _23740_/D VGND VGND VPWR VPWR _19398_/A sky130_fd_sc_hd__dfxtp_4
X_20952_ _24229_/Q _14620_/A _15915_/B _24771_/Q _15685_/X VGND VGND VPWR VPWR _20952_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__16399__B1 _16398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ _23689_/CLK _19603_/X VGND VGND VPWR VPWR _23671_/Q sky130_fd_sc_hd__dfxtp_4
X_20883_ _20900_/A VGND VGND VPWR VPWR _20889_/B sky130_fd_sc_hd__buf_2
XFILLER_53_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19337__B1 _19291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11770__A _25530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25410_ _25020_/CLK _25410_/D HRESETn VGND VGND VPWR VPWR _25410_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22622_ _22736_/A _22619_/X _22622_/C VGND VGND VPWR VPWR _22622_/X sky130_fd_sc_hd__and3_4
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21695__A1 _21512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25341_ _24868_/CLK _25341_/D HRESETn VGND VGND VPWR VPWR _12314_/A sky130_fd_sc_hd__dfrtp_4
X_22553_ _24609_/Q _22592_/B VGND VGND VPWR VPWR _22553_/X sky130_fd_sc_hd__or2_4
XANTENNA__21695__B2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21504_ _21504_/A _21504_/B VGND VGND VPWR VPWR _21504_/X sky130_fd_sc_hd__and2_4
XFILLER_107_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25272_ _25508_/CLK _25272_/D HRESETn VGND VGND VPWR VPWR _11656_/A sky130_fd_sc_hd__dfrtp_4
X_22484_ _22484_/A _22644_/B VGND VGND VPWR VPWR _22484_/X sky130_fd_sc_hd__or2_4
XANTENNA__16571__B1 _16401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25393__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24223_ _24715_/CLK _24223_/D HRESETn VGND VGND VPWR VPWR _24223_/Q sky130_fd_sc_hd__dfrtp_4
X_21435_ _21280_/B _21433_/X _21296_/X _24808_/Q _22513_/B VGND VGND VPWR VPWR _21435_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16073__A _24704_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25322__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24154_ _24643_/CLK _24154_/D HRESETn VGND VGND VPWR VPWR _18416_/A sky130_fd_sc_hd__dfrtp_4
X_21366_ _21366_/A _21498_/A VGND VGND VPWR VPWR _21366_/X sky130_fd_sc_hd__and2_4
XFILLER_68_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23105_ _21303_/X VGND VGND VPWR VPWR _23105_/X sky130_fd_sc_hd__buf_2
X_20317_ _18237_/A VGND VGND VPWR VPWR _20317_/X sky130_fd_sc_hd__buf_2
X_24085_ _25301_/CLK _24085_/D HRESETn VGND VGND VPWR VPWR _11991_/A sky130_fd_sc_hd__dfrtp_4
X_21297_ _21314_/A VGND VGND VPWR VPWR _22747_/B sky130_fd_sc_hd__buf_2
XANTENNA__22947__A1 _21409_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21419__A _21418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23036_ _24795_/Q _23101_/B VGND VGND VPWR VPWR _23036_/X sky130_fd_sc_hd__or2_4
X_20248_ _20247_/Y _20245_/X _18267_/X _20245_/X VGND VGND VPWR VPWR _23438_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22411__A3 _22396_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16626__A1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20179_ _20179_/A VGND VGND VPWR VPWR _21765_/B sky130_fd_sc_hd__inv_2
XFILLER_76_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_8_0_HCLK_A clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_21_0_HCLK clkbuf_8_21_0_HCLK/A VGND VGND VPWR VPWR _25199_/CLK sky130_fd_sc_hd__clkbuf_1
X_24987_ _24995_/CLK _15343_/X HRESETn VGND VGND VPWR VPWR _24987_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18728__A _18675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_84_0_HCLK clkbuf_7_42_0_HCLK/X VGND VGND VPWR VPWR _24955_/CLK sky130_fd_sc_hd__clkbuf_1
X_14740_ _22038_/A _14740_/B VGND VGND VPWR VPWR _14740_/X sky130_fd_sc_hd__or2_4
XANTENNA__24275__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11952_ _19629_/A VGND VGND VPWR VPWR _11952_/X sky130_fd_sc_hd__buf_2
XFILLER_57_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23938_ _24364_/CLK _20569_/Y HRESETn VGND VGND VPWR VPWR _20566_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24204__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14671_ _14670_/X VGND VGND VPWR VPWR _14671_/X sky130_fd_sc_hd__buf_2
X_11883_ _11878_/A VGND VGND VPWR VPWR _11883_/Y sky130_fd_sc_hd__inv_2
X_23869_ _23869_/CLK _19035_/X VGND VGND VPWR VPWR _23869_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19328__B1 _19191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16410_ HWDATA[17] VGND VGND VPWR VPWR _16410_/X sky130_fd_sc_hd__buf_2
XFILLER_83_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13622_ _18057_/A _13621_/X _18057_/A _13621_/X VGND VGND VPWR VPWR _13623_/A sky130_fd_sc_hd__a2bb2o_4
X_17390_ _20620_/A _20620_/B VGND VGND VPWR VPWR _20621_/A sky130_fd_sc_hd__or2_4
XFILLER_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16341_ _16339_/Y _16337_/X _16340_/X _16337_/X VGND VGND VPWR VPWR _16341_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13553_ _13551_/Y _25076_/Q _13846_/A _14560_/A VGND VGND VPWR VPWR _13553_/X sky130_fd_sc_hd__a2bb2o_4
X_25539_ _23384_/CLK _11705_/X HRESETn VGND VGND VPWR VPWR _25539_/Q sky130_fd_sc_hd__dfrtp_4
X_12504_ _12280_/Y _12509_/B VGND VGND VPWR VPWR _12505_/C sky130_fd_sc_hd__nand2_4
X_19060_ _23860_/Q VGND VGND VPWR VPWR _19060_/Y sky130_fd_sc_hd__inv_2
X_16272_ _15646_/X _15993_/Y _16270_/X _21003_/A _16271_/X VGND VGND VPWR VPWR _16272_/X
+ sky130_fd_sc_hd__a32o_4
X_13484_ _13484_/A VGND VGND VPWR VPWR _13484_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15223_ _15219_/B _15223_/B VGND VGND VPWR VPWR _15228_/B sky130_fd_sc_hd__or2_4
X_18011_ _18215_/A _19157_/A VGND VGND VPWR VPWR _18012_/C sky130_fd_sc_hd__or2_4
X_12435_ _12284_/A _12434_/Y VGND VGND VPWR VPWR _12435_/X sky130_fd_sc_hd__or2_4
XANTENNA__25063__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15154_ _15153_/Y _24570_/Q _15422_/A _15125_/Y VGND VGND VPWR VPWR _15154_/X sky130_fd_sc_hd__a2bb2o_4
X_12366_ _24827_/Q VGND VGND VPWR VPWR _12366_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16314__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14105_ _25212_/Q VGND VGND VPWR VPWR _14106_/C sky130_fd_sc_hd__inv_2
XANTENNA__19294__A _18996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20661__A2 _17404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15085_ _15365_/A _24583_/Q _15083_/Y _24583_/Q VGND VGND VPWR VPWR _15085_/X sky130_fd_sc_hd__a2bb2o_4
X_19962_ _21795_/B _19957_/X _19625_/X _19957_/X VGND VGND VPWR VPWR _23544_/D sky130_fd_sc_hd__a2bb2o_4
X_12297_ _25349_/Q VGND VGND VPWR VPWR _13023_/A sky130_fd_sc_hd__inv_2
X_14036_ _14036_/A _14070_/B _14036_/C VGND VGND VPWR VPWR _14543_/C sky130_fd_sc_hd__or3_4
X_18913_ _23911_/Q VGND VGND VPWR VPWR _18913_/Y sky130_fd_sc_hd__inv_2
X_19893_ _19892_/Y _19890_/X _19615_/X _19890_/X VGND VGND VPWR VPWR _23571_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20233__A _20232_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23247__C _22812_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11855__A _25509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18844_ _18828_/X _18833_/X _18838_/X _18843_/X VGND VGND VPWR VPWR _18844_/X sky130_fd_sc_hd__or4_4
XFILLER_67_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21048__B _21048_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18775_ _24126_/Q _18774_/Y VGND VGND VPWR VPWR _18775_/X sky130_fd_sc_hd__or2_4
XFILLER_62_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15987_ _12224_/Y _15982_/X _15986_/X _15982_/X VGND VGND VPWR VPWR _15987_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17726_ _17722_/X _17725_/X _17722_/X _17725_/X VGND VGND VPWR VPWR _17726_/X sky130_fd_sc_hd__a2bb2o_4
X_14938_ _24997_/Q _24403_/Q _15278_/A _14937_/Y VGND VGND VPWR VPWR _14938_/X sky130_fd_sc_hd__o22a_4
XFILLER_110_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17261__B _17261_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17657_ _17580_/A _17657_/B VGND VGND VPWR VPWR _17658_/C sky130_fd_sc_hd__or2_4
X_14869_ _14869_/A VGND VGND VPWR VPWR _14869_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19319__B1 _19294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16608_ _16608_/A VGND VGND VPWR VPWR _16608_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17588_ _17617_/A _17588_/B _17588_/C VGND VGND VPWR VPWR _17588_/X sky130_fd_sc_hd__and3_4
XFILLER_35_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23998__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19327_ _23766_/Q VGND VGND VPWR VPWR _19327_/Y sky130_fd_sc_hd__inv_2
X_16539_ _24534_/Q VGND VGND VPWR VPWR _16539_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19258_ _19258_/A VGND VGND VPWR VPWR _21373_/B sky130_fd_sc_hd__inv_2
XANTENNA__23482__CLK _23498_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21429__A1 _16640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18209_ _18177_/A _18205_/X _18209_/C VGND VGND VPWR VPWR _18209_/X sky130_fd_sc_hd__or3_4
XFILLER_129_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21429__B2 _21428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19189_ _19187_/Y _19188_/X _19077_/X _19188_/X VGND VGND VPWR VPWR _23815_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14406__A _14406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13310__A _13310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21220_ _21220_/A _21220_/B _21220_/C VGND VGND VPWR VPWR _21220_/X sky130_fd_sc_hd__and3_4
XFILLER_30_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22623__A _22623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21151_ _16539_/Y _15852_/Y _21314_/A _21150_/X VGND VGND VPWR VPWR _21151_/X sky130_fd_sc_hd__a211o_4
XANTENNA__14208__A1_N _14207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17717__A _17717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20102_ _21256_/B _20095_/X _19841_/X _20095_/A VGND VGND VPWR VPWR _23493_/D sky130_fd_sc_hd__a2bb2o_4
X_21082_ _24807_/Q _21067_/X _21024_/X _21081_/X VGND VGND VPWR VPWR _21082_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24786__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20033_ _20033_/A VGND VGND VPWR VPWR _21789_/B sky130_fd_sc_hd__inv_2
XFILLER_119_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24910_ _24025_/CLK _24910_/D HRESETn VGND VGND VPWR VPWR _15559_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_112_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24715__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_1_0_HCLK_A clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24841_ _24840_/CLK _15776_/X HRESETn VGND VGND VPWR VPWR _24841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19558__B1 _19420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24772_ _24811_/CLK _24772_/D HRESETn VGND VGND VPWR VPWR _24772_/Q sky130_fd_sc_hd__dfrtp_4
X_21984_ _21984_/A _21862_/X _21875_/X _21983_/Y VGND VGND VPWR VPWR HRDATA[4] sky130_fd_sc_hd__or4_4
XFILLER_39_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23723_ _23869_/CLK _19450_/X VGND VGND VPWR VPWR _17989_/B sky130_fd_sc_hd__dfxtp_4
X_20935_ _24056_/Q _20931_/X _20939_/B VGND VGND VPWR VPWR _20935_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_57_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ _24197_/CLK _19656_/X VGND VGND VPWR VPWR _23654_/Q sky130_fd_sc_hd__dfxtp_4
X_20866_ _20860_/X _20862_/Y _24476_/Q _20865_/X VGND VGND VPWR VPWR _24039_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22605_ _22589_/Y _22594_/Y _22602_/Y _21437_/X _22604_/X VGND VGND VPWR VPWR _22606_/A
+ sky130_fd_sc_hd__a32o_4
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23585_ _23581_/CLK _19855_/X VGND VGND VPWR VPWR _19854_/A sky130_fd_sc_hd__dfxtp_4
X_20797_ _15570_/Y _20676_/X _20770_/A _20796_/Y VGND VGND VPWR VPWR _20797_/X sky130_fd_sc_hd__o22a_4
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25503__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22517__B _22782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25324_ _24836_/CLK _25324_/D HRESETn VGND VGND VPWR VPWR _25324_/Q sky130_fd_sc_hd__dfrtp_4
X_22536_ _17350_/C _22534_/X _22535_/Y VGND VGND VPWR VPWR _22536_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21421__B _21420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25255_ _25255_/CLK _13826_/X HRESETn VGND VGND VPWR VPWR _25255_/Q sky130_fd_sc_hd__dfrtp_4
X_22467_ _21066_/A VGND VGND VPWR VPWR _22467_/X sky130_fd_sc_hd__buf_2
XANTENNA__11908__A1 _13678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12220_ _12220_/A VGND VGND VPWR VPWR _12220_/X sky130_fd_sc_hd__buf_2
X_24206_ _24290_/CLK _18284_/X HRESETn VGND VGND VPWR VPWR _17729_/A sky130_fd_sc_hd__dfrtp_4
X_21418_ _22598_/B VGND VGND VPWR VPWR _21418_/X sky130_fd_sc_hd__buf_2
XANTENNA__18297__B1 _21491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18836__A2 _24121_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25186_ _24942_/CLK _14230_/X HRESETn VGND VGND VPWR VPWR _25186_/Q sky130_fd_sc_hd__dfstp_4
X_22398_ _24252_/Q _21095_/X _23314_/B VGND VGND VPWR VPWR _22398_/X sky130_fd_sc_hd__o21a_4
XFILLER_118_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12151_ _12151_/A _12148_/A VGND VGND VPWR VPWR _12153_/A sky130_fd_sc_hd__and2_4
XFILLER_120_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24137_ _24136_/CLK _24137_/D HRESETn VGND VGND VPWR VPWR _24137_/Q sky130_fd_sc_hd__dfrtp_4
X_21349_ _21348_/X VGND VGND VPWR VPWR _21349_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21149__A _16622_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12082_ _12081_/Y _12079_/X _11847_/X _12079_/X VGND VGND VPWR VPWR _12082_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17346__B _17346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24068_ _24069_/CLK _20520_/X HRESETn VGND VGND VPWR VPWR _24068_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13530__B1 SCLK_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15910_ _15705_/X _15894_/X _15845_/X _24772_/Q _15864_/A VGND VGND VPWR VPWR _24772_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_78_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24456__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23019_ _24455_/Q _23019_/B _23019_/C VGND VGND VPWR VPWR _23019_/X sky130_fd_sc_hd__and3_4
X_16890_ _16137_/Y _17744_/A _16137_/Y _17744_/A VGND VGND VPWR VPWR _16890_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13593__C _11714_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17272__A1 _17235_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23364__A _21007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15841_ _12344_/Y _15833_/X _15840_/X _15809_/A VGND VGND VPWR VPWR _24808_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18458__A _24168_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23345__A1 _11970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18560_ _18475_/B _18559_/X VGND VGND VPWR VPWR _18580_/A sky130_fd_sc_hd__or2_4
XANTENNA__23083__B _23019_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12984_ _13043_/A VGND VGND VPWR VPWR _13002_/B sky130_fd_sc_hd__buf_2
X_15772_ _15749_/X _15765_/X _15647_/X _24842_/Q _15711_/A VGND VGND VPWR VPWR _15772_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_45_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17511_ _25531_/Q _24302_/Q _11766_/Y _17616_/A VGND VGND VPWR VPWR _17514_/C sky130_fd_sc_hd__o22a_4
X_11935_ _11947_/A VGND VGND VPWR VPWR _11935_/X sky130_fd_sc_hd__buf_2
X_14723_ _14722_/X VGND VGND VPWR VPWR _14723_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18491_ _18456_/X _18503_/B VGND VGND VPWR VPWR _18491_/X sky130_fd_sc_hd__or2_4
XFILLER_45_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14654_ _13605_/B _14638_/X _14648_/X _14653_/X VGND VGND VPWR VPWR _25063_/D sky130_fd_sc_hd__a22oi_4
X_17442_ _11865_/X VGND VGND VPWR VPWR _17442_/X sky130_fd_sc_hd__buf_2
X_11866_ _11865_/X VGND VGND VPWR VPWR _11867_/A sky130_fd_sc_hd__buf_2
XANTENNA__22708__A _22708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13605_ _14785_/A _13605_/B VGND VGND VPWR VPWR _13605_/X sky130_fd_sc_hd__and2_4
XFILLER_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21612__A _21612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14585_ _14581_/B _14557_/X _14584_/X _13770_/X _14558_/X VGND VGND VPWR VPWR _14585_/X
+ sky130_fd_sc_hd__a32o_4
X_17373_ _17370_/A _17369_/B _17373_/C VGND VGND VPWR VPWR _17373_/X sky130_fd_sc_hd__and3_4
XFILLER_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11797_ _11793_/Y _11795_/X _11796_/X _11795_/X VGND VGND VPWR VPWR _25523_/D sky130_fd_sc_hd__a2bb2o_4
X_19112_ _19106_/Y VGND VGND VPWR VPWR _19112_/X sky130_fd_sc_hd__buf_2
XANTENNA__25244__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13536_ _13536_/A VGND VGND VPWR VPWR _13536_/Y sky130_fd_sc_hd__inv_2
X_16324_ _16324_/A VGND VGND VPWR VPWR _16324_/X sky130_fd_sc_hd__buf_2
XFILLER_9_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16255_ _16253_/Y _16254_/X _16061_/X _16254_/X VGND VGND VPWR VPWR _16255_/X sky130_fd_sc_hd__a2bb2o_4
X_19043_ _19042_/Y _19040_/X _18993_/X _19040_/X VGND VGND VPWR VPWR _19043_/X sky130_fd_sc_hd__a2bb2o_4
X_13467_ _12050_/A _15991_/B _11716_/A _13593_/D VGND VGND VPWR VPWR _13467_/X sky130_fd_sc_hd__or4_4
XFILLER_51_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18921__A _23908_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15206_ _15199_/A _15203_/B _15205_/X VGND VGND VPWR VPWR _15207_/A sky130_fd_sc_hd__or3_4
X_12418_ _12184_/A _12417_/Y VGND VGND VPWR VPWR _12420_/B sky130_fd_sc_hd__or2_4
X_16186_ _16192_/A VGND VGND VPWR VPWR _16187_/A sky130_fd_sc_hd__buf_2
XFILLER_103_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13398_ _13177_/Y _13398_/B _13398_/C VGND VGND VPWR VPWR _13398_/X sky130_fd_sc_hd__and3_4
XFILLER_138_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15137_ _24980_/Q VGND VGND VPWR VPWR _15369_/A sky130_fd_sc_hd__inv_2
X_12349_ _12349_/A VGND VGND VPWR VPWR _12349_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16441__A HWDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15068_ _15068_/A _14947_/Y _15068_/C _15211_/A VGND VGND VPWR VPWR _15068_/X sky130_fd_sc_hd__or4_4
X_19945_ _19945_/A VGND VGND VPWR VPWR _19945_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13784__B _16725_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14019_ _13982_/A _13983_/X _13977_/X _13980_/Y VGND VGND VPWR VPWR _14020_/B sky130_fd_sc_hd__or4_4
XANTENNA__19788__B1 _19787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24197__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19876_ _19875_/Y _19873_/X _19622_/X _19873_/X VGND VGND VPWR VPWR _19876_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24126__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18827_ _16469_/Y _24141_/Q _16469_/Y _24141_/Q VGND VGND VPWR VPWR _18827_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18758_ _18758_/A _18758_/B VGND VGND VPWR VPWR _18758_/Y sky130_fd_sc_hd__nand2_4
XFILLER_110_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17709_ _17713_/A VGND VGND VPWR VPWR _17709_/Y sky130_fd_sc_hd__inv_2
X_18689_ _18768_/A _18765_/A _18610_/Y _18656_/Y VGND VGND VPWR VPWR _18692_/C sky130_fd_sc_hd__or4_4
X_20720_ _20719_/X VGND VGND VPWR VPWR _20720_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16774__B1 _16600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20651_ _17398_/B _20650_/Y _20651_/C VGND VGND VPWR VPWR _20651_/X sky130_fd_sc_hd__and3_4
XANTENNA__22847__B1 _11790_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23370_ _23370_/CLK HSEL VGND VGND VPWR VPWR _23333_/B sky130_fd_sc_hd__dfxtp_4
X_20582_ _14416_/A _20582_/B VGND VGND VPWR VPWR _20582_/X sky130_fd_sc_hd__or2_4
XFILLER_17_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16526__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22321_ _22320_/Y _21336_/A _14218_/Y _14221_/A VGND VGND VPWR VPWR _22321_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13040__A _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25040_ _25043_/CLK _25040_/D HRESETn VGND VGND VPWR VPWR _14817_/C sky130_fd_sc_hd__dfrtp_4
X_22252_ _18293_/B _19870_/Y VGND VGND VPWR VPWR _22254_/B sky130_fd_sc_hd__or2_4
XFILLER_129_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24967__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22353__A _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21203_ _13817_/A _21202_/Y _24213_/Q _13817_/A VGND VGND VPWR VPWR _21203_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21822__A1 _21815_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22183_ _22183_/A _21293_/A VGND VGND VPWR VPWR _22183_/X sky130_fd_sc_hd__or2_4
X_21134_ _13789_/B _24178_/Q _23344_/B _12059_/X VGND VGND VPWR VPWR _21135_/B sky130_fd_sc_hd__o22a_4
XFILLER_63_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21065_ _21065_/A _21017_/B VGND VGND VPWR VPWR _21065_/X sky130_fd_sc_hd__or2_4
XFILLER_119_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20016_ _23526_/Q VGND VGND VPWR VPWR _20016_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24824_ _24852_/CLK _24824_/D HRESETn VGND VGND VPWR VPWR _24824_/Q sky130_fd_sc_hd__dfrtp_4
X_24755_ _24759_/CLK _24755_/D HRESETn VGND VGND VPWR VPWR _12257_/A sky130_fd_sc_hd__dfrtp_4
X_21967_ _21967_/A _13815_/X VGND VGND VPWR VPWR _21967_/X sky130_fd_sc_hd__or2_4
XFILLER_55_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _16371_/A _11720_/B VGND VGND VPWR VPWR _16079_/A sky130_fd_sc_hd__or2_4
XFILLER_76_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13215__A _13457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23706_ _23682_/CLK _23706_/D VGND VGND VPWR VPWR _23706_/Q sky130_fd_sc_hd__dfxtp_4
X_20918_ _13664_/A VGND VGND VPWR VPWR _20918_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16765__B1 _15745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24686_ _24689_/CLK _16121_/X HRESETn VGND VGND VPWR VPWR _22865_/A sky130_fd_sc_hd__dfrtp_4
X_21898_ _14693_/A _21896_/X _21897_/X VGND VGND VPWR VPWR _21898_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_158_0_HCLK clkbuf_7_79_0_HCLK/X VGND VGND VPWR VPWR _24267_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _17445_/B VGND VGND VPWR VPWR _11970_/C sky130_fd_sc_hd__buf_2
XPHY_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23637_ _24186_/CLK _23637_/D VGND VGND VPWR VPWR _19702_/A sky130_fd_sc_hd__dfxtp_4
X_20849_ _16702_/Y _20836_/X _20845_/X _20848_/X VGND VGND VPWR VPWR _20850_/A sky130_fd_sc_hd__o22a_4
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ _25142_/Q _14348_/Y _25141_/Q _14344_/X VGND VGND VPWR VPWR _14370_/X sky130_fd_sc_hd__o22a_4
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16517__B1 _16143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23568_ _23533_/CLK _23568_/D VGND VGND VPWR VPWR _23568_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _13421_/A _13319_/X _13320_/X VGND VGND VPWR VPWR _13321_/X sky130_fd_sc_hd__and3_4
X_25307_ _25305_/CLK _25307_/D HRESETn VGND VGND VPWR VPWR _25307_/Q sky130_fd_sc_hd__dfrtp_4
X_22519_ _22488_/X _22492_/X _22498_/Y _22518_/X VGND VGND VPWR VPWR HRDATA[9] sky130_fd_sc_hd__a211o_4
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23499_ _23498_/CLK _23499_/D VGND VGND VPWR VPWR _23499_/Q sky130_fd_sc_hd__dfxtp_4
X_16040_ _16060_/A VGND VGND VPWR VPWR _16040_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13252_ _13248_/A VGND VGND VPWR VPWR _13395_/A sky130_fd_sc_hd__buf_2
X_25238_ _25192_/CLK _13868_/X HRESETn VGND VGND VPWR VPWR _20663_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23263__B1 _12546_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23359__A _21002_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22263__A _22263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18460__B _18460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12203_ _12282_/B VGND VGND VPWR VPWR _12203_/X sky130_fd_sc_hd__buf_2
X_13183_ _13180_/A _13183_/B VGND VGND VPWR VPWR _13183_/X sky130_fd_sc_hd__or2_4
XANTENNA__24637__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25169_ _25461_/CLK _25169_/D HRESETn VGND VGND VPWR VPWR _13522_/D sky130_fd_sc_hd__dfrtp_4
X_12134_ _12134_/A VGND VGND VPWR VPWR _12134_/Y sky130_fd_sc_hd__inv_2
X_17991_ _18180_/A _23891_/Q VGND VGND VPWR VPWR _17992_/C sky130_fd_sc_hd__or2_4
X_19730_ _19729_/Y VGND VGND VPWR VPWR _19730_/X sky130_fd_sc_hd__buf_2
XFILLER_81_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24290__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12065_ _16453_/A VGND VGND VPWR VPWR _21559_/A sky130_fd_sc_hd__buf_2
X_16942_ _16100_/Y _17740_/A _16115_/A _16941_/Y VGND VGND VPWR VPWR _16942_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21577__B1 _22444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23094__A _23071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19661_ _19683_/A _19683_/B _18922_/X VGND VGND VPWR VPWR _19661_/X sky130_fd_sc_hd__or3_4
XFILLER_77_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21041__A2 _21021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16873_ _16871_/Y _16868_/X _16872_/X _16868_/X VGND VGND VPWR VPWR _16873_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18612_ _18719_/A VGND VGND VPWR VPWR _18696_/A sky130_fd_sc_hd__inv_2
X_15824_ _22873_/B VGND VGND VPWR VPWR _15824_/X sky130_fd_sc_hd__buf_2
XANTENNA__15605__A _15588_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19592_ _21963_/C VGND VGND VPWR VPWR _22046_/A sky130_fd_sc_hd__inv_2
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25496__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18543_ _18541_/A _18540_/B _18542_/Y VGND VGND VPWR VPWR _24161_/D sky130_fd_sc_hd__and3_4
Xclkbuf_7_54_0_HCLK clkbuf_7_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12967_ _12964_/A _12960_/B _12967_/C VGND VGND VPWR VPWR _12967_/X sky130_fd_sc_hd__and3_4
X_15755_ _12523_/Y _15754_/X _11822_/X _15754_/X VGND VGND VPWR VPWR _15755_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22541__A2 _22422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25425__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11918_ _25499_/Q _11916_/X _11910_/X _11917_/Y VGND VGND VPWR VPWR _11918_/X sky130_fd_sc_hd__o22a_4
X_14706_ _14705_/X VGND VGND VPWR VPWR _14707_/A sky130_fd_sc_hd__buf_2
X_18474_ _24145_/Q VGND VGND VPWR VPWR _18475_/D sky130_fd_sc_hd__inv_2
X_12898_ _12852_/X _12862_/X _12886_/A VGND VGND VPWR VPWR _12898_/X sky130_fd_sc_hd__o21a_4
X_15686_ _24771_/Q _15683_/Y _15685_/X _13591_/Y VGND VGND VPWR VPWR _15687_/C sky130_fd_sc_hd__a211o_4
XANTENNA__16756__B1 _16408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17425_ _17432_/A VGND VGND VPWR VPWR _17425_/X sky130_fd_sc_hd__buf_2
XANTENNA__16236__A1_N _16234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11849_ _11844_/Y _11836_/X _11847_/X _11848_/X VGND VGND VPWR VPWR _11849_/X sky130_fd_sc_hd__a2bb2o_4
X_14637_ _18057_/A VGND VGND VPWR VPWR _17957_/A sky130_fd_sc_hd__buf_2
XFILLER_18_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14568_ _14592_/A _14592_/B VGND VGND VPWR VPWR _14569_/A sky130_fd_sc_hd__or2_4
X_17356_ _17350_/C _17355_/X _17289_/A _17352_/B VGND VGND VPWR VPWR _17357_/A sky130_fd_sc_hd__a211o_4
XANTENNA__13779__B _14219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15492__A1_N _11707_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16307_ _16305_/Y _16303_/X _16306_/X _16303_/X VGND VGND VPWR VPWR _24622_/D sky130_fd_sc_hd__a2bb2o_4
X_13519_ _12026_/X VGND VGND VPWR VPWR _20958_/B sky130_fd_sc_hd__buf_2
X_14499_ _23379_/Q _20459_/B _14497_/X _23919_/D _14498_/Y VGND VGND VPWR VPWR _14499_/X
+ sky130_fd_sc_hd__a32o_4
X_17287_ _17279_/A VGND VGND VPWR VPWR _17289_/A sky130_fd_sc_hd__buf_2
XFILLER_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19026_ _19025_/Y _19023_/X _18955_/X _19023_/X VGND VGND VPWR VPWR _19026_/X sky130_fd_sc_hd__a2bb2o_4
X_16238_ _11812_/X VGND VGND VPWR VPWR _16238_/X sky130_fd_sc_hd__buf_2
XFILLER_134_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15994__B _15993_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23269__A _24765_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13795__A _16725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17267__A _17346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24378__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16169_ _16169_/A VGND VGND VPWR VPWR _16169_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24646__CLK _24581_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24307__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15495__B1 HADDR[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19928_ _19927_/Y _19923_/X _19841_/X _19923_/A VGND VGND VPWR VPWR _23557_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21517__A _23100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19859_ _19859_/A VGND VGND VPWR VPWR _19859_/X sky130_fd_sc_hd__buf_2
XFILLER_84_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22870_ _17254_/A _22424_/A _25373_/Q _22288_/X VGND VGND VPWR VPWR _22870_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16995__B1 _24708_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21821_ _21821_/A _21816_/X _21820_/X VGND VGND VPWR VPWR _21821_/X sky130_fd_sc_hd__and3_4
XFILLER_83_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23942__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24540_ _24541_/CLK _16526_/X HRESETn VGND VGND VPWR VPWR _24540_/Q sky130_fd_sc_hd__dfrtp_4
X_21752_ _21629_/A _21752_/B VGND VGND VPWR VPWR _21752_/X sky130_fd_sc_hd__or2_4
XFILLER_93_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21740__B1 _21105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20703_ _13128_/A _13128_/B _13129_/B VGND VGND VPWR VPWR _20703_/Y sky130_fd_sc_hd__a21boi_4
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24471_ _24649_/CLK _16708_/X HRESETn VGND VGND VPWR VPWR _24471_/Q sky130_fd_sc_hd__dfrtp_4
X_21683_ _20331_/A _22389_/B _23382_/Q _22390_/B VGND VGND VPWR VPWR _21683_/X sky130_fd_sc_hd__o22a_4
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23422_ _23398_/CLK _20291_/X VGND VGND VPWR VPWR _23422_/Q sky130_fd_sc_hd__dfxtp_4
X_20634_ _17403_/A VGND VGND VPWR VPWR _20651_/C sky130_fd_sc_hd__buf_2
XANTENNA__21099__A2 _21095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22296__A1 _24509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23353_ VGND VGND VPWR VPWR _23353_/HI sda_o_S5 sky130_fd_sc_hd__conb_1
X_20565_ _20565_/A VGND VGND VPWR VPWR _23937_/D sky130_fd_sc_hd__inv_2
X_22304_ _22304_/A VGND VGND VPWR VPWR _22309_/B sky130_fd_sc_hd__inv_2
X_23284_ _23282_/X _23283_/X _22132_/A VGND VGND VPWR VPWR _23284_/X sky130_fd_sc_hd__or3_4
X_20496_ _20452_/A _14063_/X _20496_/C _20496_/D VGND VGND VPWR VPWR _20496_/X sky130_fd_sc_hd__and4_4
X_25023_ _25024_/CLK _25023_/D HRESETn VGND VGND VPWR VPWR _25023_/Q sky130_fd_sc_hd__dfrtp_4
X_22235_ _22009_/A _22235_/B VGND VGND VPWR VPWR _22235_/X sky130_fd_sc_hd__or2_4
XFILLER_69_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24730__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24048__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22166_ _17369_/A _22419_/A _25426_/Q _21062_/Y VGND VGND VPWR VPWR _22166_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20074__A3 _11862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22811__A _15854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21117_ _24919_/Q _11726_/B _13771_/X _11709_/B VGND VGND VPWR VPWR _21350_/B sky130_fd_sc_hd__or4_4
X_22097_ _22097_/A VGND VGND VPWR VPWR _22097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12114__A _12119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21048_ _21048_/A _21048_/B VGND VGND VPWR VPWR _21048_/X sky130_fd_sc_hd__or2_4
XFILLER_87_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20331__A _20331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13870_ _13852_/X _13869_/X _14261_/A _13867_/X VGND VGND VPWR VPWR _13870_/X sky130_fd_sc_hd__o22a_4
X_12821_ _12819_/X _24776_/Q _25383_/Q _12820_/Y VGND VGND VPWR VPWR _12827_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24807_ _24842_/CLK _24807_/D HRESETn VGND VGND VPWR VPWR _24807_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22999_ _15025_/A _22998_/X _22885_/X VGND VGND VPWR VPWR _22999_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19924__B1 _19794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17640__A _17525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12752_ _12752_/A VGND VGND VPWR VPWR _12753_/A sky130_fd_sc_hd__inv_2
X_15540_ _24913_/Q VGND VGND VPWR VPWR _15540_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16738__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24738_ _24804_/CLK _15985_/X HRESETn VGND VGND VPWR VPWR _24738_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11650_/A _11970_/D VGND VGND VPWR VPWR _11704_/A sky130_fd_sc_hd__and2_4
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _16355_/A VGND VGND VPWR VPWR _15471_/X sky130_fd_sc_hd__buf_2
X_12683_ _12683_/A _12686_/B VGND VGND VPWR VPWR _12683_/Y sky130_fd_sc_hd__nand2_4
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24669_ _24700_/CLK _24669_/D HRESETn VGND VGND VPWR VPWR _21426_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16256__A _22089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12784__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14421_/Y _14419_/X _14391_/X _14419_/X VGND VGND VPWR VPWR _14422_/X sky130_fd_sc_hd__a2bb2o_4
X_17210_ _16329_/Y _22702_/A _16329_/Y _22702_/A VGND VGND VPWR VPWR _17211_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12379__A2_N _12296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18190_ _18046_/A _18190_/B VGND VGND VPWR VPWR _18190_/X sky130_fd_sc_hd__or2_4
XANTENNA__24889__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14353_ _14353_/A VGND VGND VPWR VPWR _14353_/Y sky130_fd_sc_hd__inv_2
X_17141_ _17143_/A _17135_/B _17141_/C VGND VGND VPWR VPWR _24369_/D sky130_fd_sc_hd__and3_4
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24818__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13304_ _13373_/A _20240_/A VGND VGND VPWR VPWR _13305_/C sky130_fd_sc_hd__or2_4
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17072_ _17025_/B _17060_/B VGND VGND VPWR VPWR _17072_/X sky130_fd_sc_hd__or2_4
X_14284_ _14283_/X VGND VGND VPWR VPWR _14284_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13235_ _13455_/A _23651_/Q VGND VGND VPWR VPWR _13238_/B sky130_fd_sc_hd__or2_4
X_16023_ _16021_/Y _16022_/X _15955_/X _16022_/X VGND VGND VPWR VPWR _16023_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13724__B1 _13714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24471__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18258__A3 _16270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21798__B1 _18299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24400__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13166_ _13190_/A _23628_/Q VGND VGND VPWR VPWR _13166_/X sky130_fd_sc_hd__or2_4
XFILLER_112_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14223__B _14223_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12117_ _12116_/Y _12114_/X _11853_/X _12114_/X VGND VGND VPWR VPWR _12117_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13097_ _13076_/A _13097_/B _13096_/Y VGND VGND VPWR VPWR _25329_/D sky130_fd_sc_hd__and3_4
X_17974_ _17973_/X _17974_/B VGND VGND VPWR VPWR _17978_/B sky130_fd_sc_hd__or2_4
XFILLER_2_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19713_ _19711_/Y _19707_/X _19645_/X _19712_/X VGND VGND VPWR VPWR _19713_/X sky130_fd_sc_hd__a2bb2o_4
X_12048_ _16183_/A VGND VGND VPWR VPWR _13533_/A sky130_fd_sc_hd__buf_2
X_16925_ _16122_/A _17758_/B _16154_/Y _24250_/Q VGND VGND VPWR VPWR _16925_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15229__B1 _15199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12959__A _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20222__B1 _19740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19644_ _23658_/Q VGND VGND VPWR VPWR _19644_/Y sky130_fd_sc_hd__inv_2
X_16856_ _16855_/Y _16796_/X _16720_/X _16796_/X VGND VGND VPWR VPWR _16856_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15807_ _15781_/X _15795_/X _15729_/X _24830_/Q _15793_/X VGND VGND VPWR VPWR _24830_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19575_ _19573_/Y _19574_/X _11952_/X _19574_/X VGND VGND VPWR VPWR _19575_/X sky130_fd_sc_hd__a2bb2o_4
X_16787_ _16786_/X VGND VGND VPWR VPWR _16787_/X sky130_fd_sc_hd__buf_2
X_13999_ _13999_/A VGND VGND VPWR VPWR _13999_/X sky130_fd_sc_hd__buf_2
XFILLER_80_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18526_ _18400_/A _18525_/Y VGND VGND VPWR VPWR _18526_/X sky130_fd_sc_hd__or2_4
XFILLER_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15738_ _12559_/Y _15735_/X _11791_/X _15735_/X VGND VGND VPWR VPWR _15738_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21722__B1 _24570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18194__A2 _18178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18457_ _24171_/Q VGND VGND VPWR VPWR _18457_/Y sky130_fd_sc_hd__inv_2
X_15669_ _15668_/X VGND VGND VPWR VPWR _15669_/X sky130_fd_sc_hd__buf_2
XANTENNA__12694__A _12565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17700__D _17447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_141_0_HCLK clkbuf_7_70_0_HCLK/X VGND VGND VPWR VPWR _23377_/CLK sky130_fd_sc_hd__clkbuf_1
X_17408_ _17387_/X _17401_/X _24323_/Q _24324_/Q _17404_/X VGND VGND VPWR VPWR _17408_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12215__B1 _12286_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18388_ _24103_/Q _18371_/A _24178_/Q _18384_/X VGND VGND VPWR VPWR _18388_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12766__A1 _25373_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17339_ _17248_/A _17338_/Y VGND VGND VPWR VPWR _17339_/X sky130_fd_sc_hd__or2_4
XANTENNA__24559__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20350_ _21792_/B _20345_/X _11948_/A _20345_/X VGND VGND VPWR VPWR _23399_/D sky130_fd_sc_hd__a2bb2o_4
X_19009_ _19009_/A VGND VGND VPWR VPWR _19009_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13715__B1 _13714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12518__B2 _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20281_ _22250_/B _20278_/X _19978_/X _20278_/X VGND VGND VPWR VPWR _23426_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14414__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22020_ _21664_/A _22020_/B VGND VGND VPWR VPWR _22022_/B sky130_fd_sc_hd__or2_4
XANTENNA__24141__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23971_ _24943_/CLK _23971_/D HRESETn VGND VGND VPWR VPWR _17389_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20213__B1 _18247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25347__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22922_ _22922_/A VGND VGND VPWR VPWR _22922_/X sky130_fd_sc_hd__buf_2
X_22853_ _22853_/A _23304_/B VGND VGND VPWR VPWR _22853_/X sky130_fd_sc_hd__or2_4
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21804_ _21670_/A _21804_/B VGND VGND VPWR VPWR _21804_/X sky130_fd_sc_hd__or2_4
XFILLER_24_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22784_ _22913_/A VGND VGND VPWR VPWR _22872_/B sky130_fd_sc_hd__buf_2
XFILLER_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19382__B2 _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24523_ _24555_/CLK _16571_/X HRESETn VGND VGND VPWR VPWR _24523_/Q sky130_fd_sc_hd__dfrtp_4
X_21735_ _16616_/Y _21570_/X _21316_/A _21734_/X VGND VGND VPWR VPWR _21735_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22269__A1 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24454_ _25024_/CLK _24454_/D HRESETn VGND VGND VPWR VPWR _15025_/A sky130_fd_sc_hd__dfrtp_4
X_21666_ _21649_/A _21664_/X _21665_/X VGND VGND VPWR VPWR _21666_/X sky130_fd_sc_hd__and3_4
XANTENNA__24982__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23405_ _24208_/CLK _23405_/D VGND VGND VPWR VPWR _20333_/A sky130_fd_sc_hd__dfxtp_4
X_20617_ _20617_/A VGND VGND VPWR VPWR _23971_/D sky130_fd_sc_hd__inv_2
XANTENNA__24911__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24385_ _24368_/CLK _24385_/D HRESETn VGND VGND VPWR VPWR _24385_/Q sky130_fd_sc_hd__dfrtp_4
X_21597_ _21622_/A VGND VGND VPWR VPWR _21630_/A sky130_fd_sc_hd__buf_2
XFILLER_138_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24229__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23336_ _23336_/A _22044_/B VGND VGND VPWR VPWR _23336_/Y sky130_fd_sc_hd__nor2_4
X_20548_ _23934_/Q _18871_/X VGND VGND VPWR VPWR _20548_/Y sky130_fd_sc_hd__nand2_4
XFILLER_137_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23267_ _23262_/Y _23266_/Y _22850_/X VGND VGND VPWR VPWR _23267_/X sky130_fd_sc_hd__o21a_4
X_20479_ _20479_/A _14207_/A _20479_/C VGND VGND VPWR VPWR _20479_/X sky130_fd_sc_hd__and3_4
X_13020_ _13002_/B _13001_/D VGND VGND VPWR VPWR _13023_/B sky130_fd_sc_hd__or2_4
X_25006_ _25001_/CLK _25006_/D HRESETn VGND VGND VPWR VPWR _14885_/A sky130_fd_sc_hd__dfrtp_4
X_22218_ _14749_/A _22214_/X _22218_/C VGND VGND VPWR VPWR _22218_/X sky130_fd_sc_hd__or3_4
XFILLER_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23198_ _13118_/A _21278_/X _24056_/Q _21302_/X VGND VGND VPWR VPWR _23199_/B sky130_fd_sc_hd__a22oi_4
X_22149_ _22035_/X _22149_/B _22149_/C _22148_/X VGND VGND VPWR VPWR HRDATA[5] sky130_fd_sc_hd__or4_4
XFILLER_126_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14971_ _14971_/A VGND VGND VPWR VPWR _14971_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16710_ _16709_/Y _16707_/X _16355_/X _16707_/X VGND VGND VPWR VPWR _24470_/D sky130_fd_sc_hd__a2bb2o_4
X_13922_ _13919_/X _13920_/X _13921_/Y VGND VGND VPWR VPWR _13930_/A sky130_fd_sc_hd__o21ai_4
X_17690_ _17662_/A _17689_/X VGND VGND VPWR VPWR _17692_/A sky130_fd_sc_hd__nand2_4
XANTENNA__25017__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16641_ _15824_/X _15643_/Y HWDATA[31] _23317_/A _16643_/A VGND VGND VPWR VPWR _16641_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_35_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13853_ _13853_/A _13851_/X VGND VGND VPWR VPWR _13853_/Y sky130_fd_sc_hd__nor2_4
XFILLER_62_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12804_ _12804_/A _12804_/B _12800_/X _12803_/X VGND VGND VPWR VPWR _12836_/A sky130_fd_sc_hd__or4_4
X_19360_ _18024_/B VGND VGND VPWR VPWR _19360_/Y sky130_fd_sc_hd__inv_2
X_16572_ _24522_/Q VGND VGND VPWR VPWR _16572_/Y sky130_fd_sc_hd__inv_2
X_13784_ _16725_/A _16725_/B _13784_/C _13784_/D VGND VGND VPWR VPWR _13784_/X sky130_fd_sc_hd__and4_4
XFILLER_43_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18311_ _17733_/A VGND VGND VPWR VPWR _18311_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15523_ _15523_/A VGND VGND VPWR VPWR _15523_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12735_ _12735_/A VGND VGND VPWR VPWR _12736_/B sky130_fd_sc_hd__inv_2
X_19291_ _19642_/A VGND VGND VPWR VPWR _19291_/X sky130_fd_sc_hd__buf_2
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18242_ _18233_/A VGND VGND VPWR VPWR _18242_/X sky130_fd_sc_hd__buf_2
XFILLER_30_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12666_ _12666_/A _12674_/B VGND VGND VPWR VPWR _12666_/X sky130_fd_sc_hd__or2_4
X_15454_ _24068_/Q _15449_/X _15441_/Y _13905_/C _15452_/X VGND VGND VPWR VPWR _15454_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_8_214_0_HCLK clkbuf_8_215_0_HCLK/A VGND VGND VPWR VPWR _24998_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19125__B2 _19106_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ _25132_/Q VGND VGND VPWR VPWR _14405_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18832__A1_N _16483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18173_ _14646_/X _18171_/X _18172_/X VGND VGND VPWR VPWR _18173_/X sky130_fd_sc_hd__and3_4
XANTENNA__24652__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _12595_/Y _12514_/A _12731_/A _24845_/Q VGND VGND VPWR VPWR _12598_/D sky130_fd_sc_hd__a2bb2o_4
X_15385_ _15128_/Y _15379_/X _15382_/B _15339_/X VGND VGND VPWR VPWR _15385_/X sky130_fd_sc_hd__a211o_4
XFILLER_106_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17136__B1 _17056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17124_ _17143_/A _17122_/X _17123_/X VGND VGND VPWR VPWR _24373_/D sky130_fd_sc_hd__and3_4
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14336_ _25153_/Q _24094_/Q _14336_/C VGND VGND VPWR VPWR _25153_/D sky130_fd_sc_hd__and3_4
XANTENNA__22680__A1 _22671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11858__A _15986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14267_ _14266_/Y _14264_/X _13797_/X _14264_/X VGND VGND VPWR VPWR _14267_/X sky130_fd_sc_hd__a2bb2o_4
X_17055_ _17020_/X VGND VGND VPWR VPWR _17384_/B sky130_fd_sc_hd__inv_2
XANTENNA__18847__A1_N _21837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13218_ _13155_/Y VGND VGND VPWR VPWR _13309_/A sky130_fd_sc_hd__buf_2
X_16006_ _16005_/Y _16003_/X _15942_/X _16003_/X VGND VGND VPWR VPWR _16006_/X sky130_fd_sc_hd__a2bb2o_4
X_14198_ _14807_/A _14210_/B VGND VGND VPWR VPWR _14200_/A sky130_fd_sc_hd__nor2_4
XANTENNA__12256__A2_N _24739_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13149_ _13186_/A _19660_/A VGND VGND VPWR VPWR _13154_/B sky130_fd_sc_hd__or2_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21067__A _21067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17957_ _17957_/A _17957_/B _17957_/C VGND VGND VPWR VPWR _17957_/X sky130_fd_sc_hd__and3_4
XFILLER_85_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15870__B1 _11749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22735__A2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25440__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16908_ _24676_/Q _24253_/Q _16146_/Y _17846_/A VGND VGND VPWR VPWR _16908_/X sky130_fd_sc_hd__o22a_4
X_17888_ _17700_/X _17735_/B VGND VGND VPWR VPWR _17891_/A sky130_fd_sc_hd__and2_4
X_19627_ _19627_/A VGND VGND VPWR VPWR _19627_/Y sky130_fd_sc_hd__inv_2
X_16839_ _14900_/Y _16837_/X _11821_/X _16837_/X VGND VGND VPWR VPWR _24411_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25454__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19558_ _19557_/Y _19552_/X _19420_/X _19538_/X VGND VGND VPWR VPWR _23685_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22499__A1 _16246_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_24_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_24_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18509_ _18458_/Y _18508_/X VGND VGND VPWR VPWR _18517_/B sky130_fd_sc_hd__or2_4
XFILLER_0_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19489_ _19487_/Y _19483_/X _19488_/X _19470_/Y VGND VGND VPWR VPWR _19489_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14409__A _14408_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21520_ _21111_/X VGND VGND VPWR VPWR _21520_/X sky130_fd_sc_hd__buf_2
XANTENNA__13313__A _13450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22626__A _24747_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21451_ _21648_/A _20292_/Y VGND VGND VPWR VPWR _21451_/X sky130_fd_sc_hd__or2_4
XANTENNA__24393__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20402_ _23377_/Q VGND VGND VPWR VPWR _20402_/Y sky130_fd_sc_hd__inv_2
X_24170_ _24171_/CLK _18512_/X HRESETn VGND VGND VPWR VPWR _18459_/A sky130_fd_sc_hd__dfrtp_4
X_21382_ _21393_/A _21382_/B VGND VGND VPWR VPWR _21383_/C sky130_fd_sc_hd__or2_4
XANTENNA__17439__B _13789_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23121_ _22786_/A VGND VGND VPWR VPWR _23121_/X sky130_fd_sc_hd__buf_2
X_20333_ _20333_/A VGND VGND VPWR VPWR _21985_/B sky130_fd_sc_hd__inv_2
XFILLER_107_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11768__A _11777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23052_ _15579_/Y _23052_/B VGND VGND VPWR VPWR _23052_/X sky130_fd_sc_hd__and2_4
X_20264_ _21769_/B _20259_/X _19790_/A _20259_/X VGND VGND VPWR VPWR _23432_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22423__B2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22361__A _22055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22003_ _21663_/A VGND VGND VPWR VPWR _22016_/A sky130_fd_sc_hd__buf_2
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25528__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20195_ _23458_/Q VGND VGND VPWR VPWR _20195_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_106_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_213_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_23954_ _25137_/CLK _20601_/X HRESETn VGND VGND VPWR VPWR _14380_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__25110__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22905_ _22778_/A _22905_/B _22905_/C _22904_/X VGND VGND VPWR VPWR _22905_/X sky130_fd_sc_hd__or4_4
XFILLER_99_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23885_ _23869_/CLK _23885_/D VGND VGND VPWR VPWR _23885_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15613__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22836_ _24450_/Q _22836_/B _23019_/C VGND VGND VPWR VPWR _22836_/X sky130_fd_sc_hd__and3_4
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22767_ _22470_/X _22765_/X _21416_/X _24858_/Q _22766_/X VGND VGND VPWR VPWR _22768_/B
+ sky130_fd_sc_hd__a32o_4
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _12520_/A VGND VGND VPWR VPWR _12520_/Y sky130_fd_sc_hd__inv_2
X_21718_ _21718_/A VGND VGND VPWR VPWR _21718_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24506_ _24545_/CLK _16615_/X HRESETn VGND VGND VPWR VPWR _24506_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25486_ _23689_/CLK _11980_/X HRESETn VGND VGND VPWR VPWR _11653_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22698_ _16230_/A _22298_/B VGND VGND VPWR VPWR _22698_/X sky130_fd_sc_hd__or2_4
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _12451_/A VGND VGND VPWR VPWR _12451_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21440__A _15784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21649_ _21649_/A _21647_/X _21649_/C VGND VGND VPWR VPWR _21649_/X sky130_fd_sc_hd__and3_4
XFILLER_8_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24437_ _24407_/CLK _24437_/D HRESETn VGND VGND VPWR VPWR _15027_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15170_ _15198_/A _15168_/X _15170_/C VGND VGND VPWR VPWR _15170_/X sky130_fd_sc_hd__and3_4
XANTENNA__24063__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12382_ _12382_/A _12382_/B VGND VGND VPWR VPWR _12382_/X sky130_fd_sc_hd__or2_4
XFILLER_123_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24368_ _24368_/CLK _17143_/X HRESETn VGND VGND VPWR VPWR _24368_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_44_0_HCLK clkbuf_8_45_0_HCLK/A VGND VGND VPWR VPWR _25485_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_138_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14121_ _25132_/Q _14110_/X _14111_/X _14120_/Y VGND VGND VPWR VPWR _14121_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23319_ _22783_/A _23317_/Y _22786_/A _23318_/Y VGND VGND VPWR VPWR _23320_/B sky130_fd_sc_hd__o22a_4
XFILLER_67_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24299_ _25433_/CLK _24299_/D HRESETn VGND VGND VPWR VPWR _24299_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16341__B2 _16337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14052_ _14015_/X _14051_/X VGND VGND VPWR VPWR _14052_/X sky130_fd_sc_hd__or2_4
XFILLER_4_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24944__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13003_ _13005_/B VGND VGND VPWR VPWR _13004_/B sky130_fd_sc_hd__inv_2
XANTENNA__25269__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18860_ _16510_/Y _18789_/A _21837_/A _18678_/Y VGND VGND VPWR VPWR _18860_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17811_ _16941_/Y _17810_/X VGND VGND VPWR VPWR _17814_/B sky130_fd_sc_hd__or2_4
XFILLER_122_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18791_ _18799_/A _18791_/B _18791_/C VGND VGND VPWR VPWR _24124_/D sky130_fd_sc_hd__and3_4
X_17742_ _17742_/A VGND VGND VPWR VPWR _17743_/A sky130_fd_sc_hd__inv_2
XANTENNA__19043__B1 _18993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14954_ _15209_/A _16832_/A _15209_/A _16832_/A VGND VGND VPWR VPWR _14954_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13905_ _13905_/A _13905_/B _13905_/C _13904_/Y VGND VGND VPWR VPWR _13905_/X sky130_fd_sc_hd__and4_4
XFILLER_78_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17673_ _17652_/X _17673_/B _17672_/Y VGND VGND VPWR VPWR _24288_/D sky130_fd_sc_hd__and3_4
X_14885_ _14885_/A VGND VGND VPWR VPWR _14885_/Y sky130_fd_sc_hd__inv_2
X_19412_ _19412_/A VGND VGND VPWR VPWR _19412_/Y sky130_fd_sc_hd__inv_2
X_16624_ _14770_/B _16174_/B _14555_/B VGND VGND VPWR VPWR _16624_/X sky130_fd_sc_hd__o21a_4
X_13836_ _13557_/Y _13833_/X _13835_/X _13833_/X VGND VGND VPWR VPWR _13836_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19343_ _18118_/B VGND VGND VPWR VPWR _19343_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16555_ _24529_/Q VGND VGND VPWR VPWR _16555_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24833__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13767_ _20043_/C _20043_/D _20043_/C _20043_/D VGND VGND VPWR VPWR _13767_/X sky130_fd_sc_hd__a2bb2o_4
X_15506_ _15506_/A VGND VGND VPWR VPWR _15506_/Y sky130_fd_sc_hd__inv_2
X_12718_ _12706_/A _12706_/B VGND VGND VPWR VPWR _12719_/C sky130_fd_sc_hd__nand2_4
X_19274_ _21886_/B _19271_/X _16876_/X _19271_/X VGND VGND VPWR VPWR _23785_/D sky130_fd_sc_hd__a2bb2o_4
X_16486_ _16474_/A VGND VGND VPWR VPWR _16486_/X sky130_fd_sc_hd__buf_2
XANTENNA__15907__B2 _15864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13698_ _11659_/Y _13698_/B VGND VGND VPWR VPWR _13702_/B sky130_fd_sc_hd__or2_4
XANTENNA__12180__A2_N _24766_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18225_ _18097_/A _18217_/X _18224_/X VGND VGND VPWR VPWR _18225_/X sky130_fd_sc_hd__and3_4
XANTENNA__21350__A _14190_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15437_ _15449_/A VGND VGND VPWR VPWR _15437_/X sky130_fd_sc_hd__buf_2
XFILLER_54_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12649_ _12648_/X VGND VGND VPWR VPWR _25414_/D sky130_fd_sc_hd__inv_2
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18156_ _18220_/A _18154_/X _18156_/C VGND VGND VPWR VPWR _18160_/B sky130_fd_sc_hd__and3_4
XANTENNA__18857__B1 _16503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24083__D _20951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15368_ _15372_/A _15362_/X _15368_/C VGND VGND VPWR VPWR _24981_/D sky130_fd_sc_hd__and3_4
X_17107_ _17034_/A _17110_/B VGND VGND VPWR VPWR _17107_/Y sky130_fd_sc_hd__nand2_4
XFILLER_129_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14319_ _25160_/Q _14299_/Y _25159_/Q _14296_/B VGND VGND VPWR VPWR _14319_/X sky130_fd_sc_hd__o22a_4
XFILLER_32_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19755__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18087_ _18087_/A VGND VGND VPWR VPWR _18220_/A sky130_fd_sc_hd__buf_2
X_15299_ _15299_/A _15299_/B _15392_/A _15406_/A VGND VGND VPWR VPWR _15299_/X sky130_fd_sc_hd__or4_4
X_17038_ _17038_/A _17038_/B _17038_/C _16960_/Y VGND VGND VPWR VPWR _17045_/A sky130_fd_sc_hd__or4_4
XFILLER_132_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22956__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18989_ _18988_/Y VGND VGND VPWR VPWR _18989_/X sky130_fd_sc_hd__buf_2
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21525__A _21525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20951_ _25313_/Q _11650_/A _11958_/X VGND VGND VPWR VPWR _20951_/X sky130_fd_sc_hd__a21o_4
XFILLER_96_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23670_ _23689_/CLK _23670_/D VGND VGND VPWR VPWR _23670_/Q sky130_fd_sc_hd__dfxtp_4
X_20882_ _20909_/A VGND VGND VPWR VPWR _20882_/X sky130_fd_sc_hd__buf_2
XFILLER_42_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22621_ _16592_/A _21049_/X _21731_/X _22620_/X VGND VGND VPWR VPWR _22622_/C sky130_fd_sc_hd__a211o_4
XANTENNA__24574__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25340_ _24852_/CLK _25340_/D HRESETn VGND VGND VPWR VPWR _25340_/Q sky130_fd_sc_hd__dfrtp_4
X_22552_ _22476_/X _22550_/X _21285_/A _12305_/A _22551_/X VGND VGND VPWR VPWR _22552_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_50_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24503__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22356__A _14682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16020__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21503_ _13782_/X VGND VGND VPWR VPWR _21504_/B sky130_fd_sc_hd__buf_2
X_25271_ _25508_/CLK _25271_/D HRESETn VGND VGND VPWR VPWR _11669_/A sky130_fd_sc_hd__dfrtp_4
X_22483_ _22186_/A VGND VGND VPWR VPWR _22483_/X sky130_fd_sc_hd__buf_2
X_24222_ _24715_/CLK _24222_/D HRESETn VGND VGND VPWR VPWR _22507_/A sky130_fd_sc_hd__dfrtp_4
X_21434_ _23097_/A VGND VGND VPWR VPWR _22513_/B sky130_fd_sc_hd__buf_2
Xclkbuf_8_3_0_HCLK clkbuf_8_3_0_HCLK/A VGND VGND VPWR VPWR _23609_/CLK sky130_fd_sc_hd__clkbuf_1
X_24153_ _24643_/CLK _24153_/D HRESETn VGND VGND VPWR VPWR _24153_/Q sky130_fd_sc_hd__dfrtp_4
X_21365_ _21499_/B VGND VGND VPWR VPWR _21365_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17520__B1 _11855_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23104_ _23274_/A _23104_/B VGND VGND VPWR VPWR _23104_/X sky130_fd_sc_hd__and2_4
X_20316_ _21164_/B _20311_/X _20019_/X _20298_/Y VGND VGND VPWR VPWR _23412_/D sky130_fd_sc_hd__a2bb2o_4
X_24084_ _25478_/CLK _24084_/D HRESETn VGND VGND VPWR VPWR _13643_/B sky130_fd_sc_hd__dfrtp_4
X_21296_ _21295_/X VGND VGND VPWR VPWR _21296_/X sky130_fd_sc_hd__buf_2
XANTENNA__25362__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23035_ _23035_/A VGND VGND VPWR VPWR _23101_/B sky130_fd_sc_hd__buf_2
X_20247_ _23438_/Q VGND VGND VPWR VPWR _20247_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21080__B1 _21859_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20178_ _20177_/Y _20175_/X _20089_/X _20175_/X VGND VGND VPWR VPWR _23465_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15834__B1 _15627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24986_ _24995_/CLK _24986_/D HRESETn VGND VGND VPWR VPWR _24986_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11951_ _19632_/A VGND VGND VPWR VPWR _11951_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23937_ _24364_/CLK _23937_/D HRESETn VGND VGND VPWR VPWR _18875_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_72_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11882_ _25506_/Q _11869_/X _11870_/A _13678_/B VGND VGND VPWR VPWR _11882_/X sky130_fd_sc_hd__and4_4
X_14670_ _13618_/Y _13598_/X VGND VGND VPWR VPWR _14670_/X sky130_fd_sc_hd__or2_4
XANTENNA__21154__B _21154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23868_ _25485_/CLK _19041_/X VGND VGND VPWR VPWR _23868_/Q sky130_fd_sc_hd__dfxtp_4
X_13621_ _13617_/Y _13618_/Y _14661_/A VGND VGND VPWR VPWR _13621_/X sky130_fd_sc_hd__a21o_4
X_22819_ _21275_/X VGND VGND VPWR VPWR _22819_/X sky130_fd_sc_hd__buf_2
X_23799_ _23798_/CLK _19236_/X VGND VGND VPWR VPWR _13372_/B sky130_fd_sc_hd__dfxtp_4
X_16340_ HWDATA[10] VGND VGND VPWR VPWR _16340_/X sky130_fd_sc_hd__buf_2
XANTENNA__24244__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13552_ _14610_/A VGND VGND VPWR VPWR _14560_/A sky130_fd_sc_hd__inv_2
X_25538_ _24275_/CLK _11744_/X HRESETn VGND VGND VPWR VPWR _11706_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16011__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22266__A _22590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12503_ _12503_/A _12499_/X _12502_/Y VGND VGND VPWR VPWR _25422_/D sky130_fd_sc_hd__and3_4
X_13483_ _13481_/Y _13477_/X _11842_/X _13482_/X VGND VGND VPWR VPWR _25309_/D sky130_fd_sc_hd__a2bb2o_4
X_16271_ _15649_/A _16276_/B VGND VGND VPWR VPWR _16271_/X sky130_fd_sc_hd__or2_4
X_25469_ _24097_/CLK _12084_/X HRESETn VGND VGND VPWR VPWR _12083_/A sky130_fd_sc_hd__dfrtp_4
X_18010_ _18010_/A VGND VGND VPWR VPWR _18215_/A sky130_fd_sc_hd__buf_2
X_12434_ _12433_/X VGND VGND VPWR VPWR _12434_/Y sky130_fd_sc_hd__inv_2
X_15222_ _15219_/C _15211_/B VGND VGND VPWR VPWR _15223_/B sky130_fd_sc_hd__or2_4
XANTENNA__16589__A1_N _16587_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18839__B1 _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12365_ _12363_/Y _24811_/Q _25350_/Q _12364_/Y VGND VGND VPWR VPWR _12365_/X sky130_fd_sc_hd__a2bb2o_4
X_15153_ _24966_/Q VGND VGND VPWR VPWR _15153_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17511__B1 _11766_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14104_ _14103_/X VGND VGND VPWR VPWR _14106_/B sky130_fd_sc_hd__inv_2
XFILLER_4_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15084_ _15083_/Y VGND VGND VPWR VPWR _15365_/A sky130_fd_sc_hd__buf_2
X_19961_ _23544_/Q VGND VGND VPWR VPWR _21795_/B sky130_fd_sc_hd__inv_2
XANTENNA__23097__A _23097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12296_ _12296_/A VGND VGND VPWR VPWR _12296_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22399__B1 _22397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14035_ _14035_/A VGND VGND VPWR VPWR _14036_/C sky130_fd_sc_hd__inv_2
X_18912_ _21755_/B _18907_/X _16881_/X _18907_/X VGND VGND VPWR VPWR _18912_/X sky130_fd_sc_hd__a2bb2o_4
X_19892_ _23571_/Q VGND VGND VPWR VPWR _19892_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25032__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18843_ _18839_/X _18843_/B _18843_/C _18842_/X VGND VGND VPWR VPWR _18843_/X sky130_fd_sc_hd__or4_4
XFILLER_67_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15825__B1 _24818_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18774_ _18774_/A VGND VGND VPWR VPWR _18774_/Y sky130_fd_sc_hd__inv_2
X_15986_ _15986_/A VGND VGND VPWR VPWR _15986_/X sky130_fd_sc_hd__buf_2
XFILLER_48_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17725_ _24205_/Q _17710_/X _17724_/Y VGND VGND VPWR VPWR _17725_/X sky130_fd_sc_hd__o21a_4
X_14937_ _24403_/Q VGND VGND VPWR VPWR _14937_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16439__A _24570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17656_ _24291_/Q _17656_/B VGND VGND VPWR VPWR _17656_/X sky130_fd_sc_hd__or2_4
X_14868_ _24940_/Q VGND VGND VPWR VPWR _14868_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17261__C _17235_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16250__B1 _16147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16607_ _16606_/Y _16601_/X _16521_/X _16601_/X VGND VGND VPWR VPWR _16607_/X sky130_fd_sc_hd__a2bb2o_4
X_13819_ _13771_/X _24065_/Q _13774_/Y _18235_/A VGND VGND VPWR VPWR _13820_/A sky130_fd_sc_hd__and4_4
X_17587_ _24309_/Q _17586_/B VGND VGND VPWR VPWR _17588_/C sky130_fd_sc_hd__nand2_4
XANTENNA__21126__A1 _21350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14799_ _14813_/C _14798_/X _14799_/C VGND VGND VPWR VPWR _14799_/X sky130_fd_sc_hd__or3_4
X_19326_ _19324_/Y _19325_/X _19212_/X _19325_/X VGND VGND VPWR VPWR _19326_/X sky130_fd_sc_hd__a2bb2o_4
X_16538_ _16537_/Y _16461_/A _16266_/X _16461_/A VGND VGND VPWR VPWR _24535_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12811__B1 _25376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20885__B1 _20884_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19257_ _21598_/B _19256_/X _16885_/X _19256_/X VGND VGND VPWR VPWR _19257_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22607__C _22586_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16469_ _16469_/A VGND VGND VPWR VPWR _16469_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17179__A2_N _17252_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16174__A _14555_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18208_ _18176_/A _18208_/B _18208_/C VGND VGND VPWR VPWR _18209_/C sky130_fd_sc_hd__and3_4
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13367__B2 _11965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19188_ _19175_/Y VGND VGND VPWR VPWR _19188_/X sky130_fd_sc_hd__buf_2
XANTENNA__14406__B _18895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18139_ _18024_/A _18139_/B VGND VGND VPWR VPWR _18139_/X sky130_fd_sc_hd__or2_4
XFILLER_89_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22910__A1_N _17254_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21150_ _16448_/A _15852_/A _21314_/B VGND VGND VPWR VPWR _21150_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_90_0_HCLK clkbuf_8_91_0_HCLK/A VGND VGND VPWR VPWR _24171_/CLK sky130_fd_sc_hd__clkbuf_1
X_20101_ _20101_/A VGND VGND VPWR VPWR _21256_/B sky130_fd_sc_hd__inv_2
X_21081_ _23069_/B _21073_/X _21080_/X VGND VGND VPWR VPWR _21081_/X sky130_fd_sc_hd__and3_4
XFILLER_99_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20032_ _21920_/B _20029_/X _19985_/X _20029_/X VGND VGND VPWR VPWR _23521_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24840_ _24840_/CLK _15778_/X HRESETn VGND VGND VPWR VPWR _20674_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21983_ _21982_/X VGND VGND VPWR VPWR _21983_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24755__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24771_ _23805_/CLK _15921_/X HRESETn VGND VGND VPWR VPWR _24771_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12877__A _12602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16349__A _22273_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11781__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20934_ _13666_/X VGND VGND VPWR VPWR _20939_/B sky130_fd_sc_hd__inv_2
XFILLER_96_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23722_ _23722_/CLK _23722_/D VGND VGND VPWR VPWR _18036_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ _20864_/X VGND VGND VPWR VPWR _20865_/X sky130_fd_sc_hd__buf_2
XFILLER_54_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13055__B1 _13031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23653_ _24197_/CLK _19659_/X VGND VGND VPWR VPWR _19657_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22604_ _12842_/A _22565_/X _22603_/X VGND VGND VPWR VPWR _22604_/X sky130_fd_sc_hd__o21a_4
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23584_ _23581_/CLK _19857_/X VGND VGND VPWR VPWR _23584_/Q sky130_fd_sc_hd__dfxtp_4
X_20796_ _13118_/A _20792_/X _20800_/B VGND VGND VPWR VPWR _20796_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_126_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22535_ _24039_/Q _21302_/A _24007_/Q _21304_/X VGND VGND VPWR VPWR _22535_/Y sky130_fd_sc_hd__a22oi_4
X_25323_ _25351_/CLK _25323_/D HRESETn VGND VGND VPWR VPWR _25323_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15347__A2 _15316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16084__A _15854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22466_ _22466_/A VGND VGND VPWR VPWR _22466_/X sky130_fd_sc_hd__buf_2
X_25254_ _25255_/CLK _13827_/X HRESETn VGND VGND VPWR VPWR _25254_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21417_ _21018_/A VGND VGND VPWR VPWR _22598_/B sky130_fd_sc_hd__buf_2
X_24205_ _24288_/CLK _18285_/X HRESETn VGND VGND VPWR VPWR _24205_/Q sky130_fd_sc_hd__dfrtp_4
X_25185_ _24942_/CLK _14232_/X HRESETn VGND VGND VPWR VPWR _14231_/A sky130_fd_sc_hd__dfstp_4
X_22397_ _11831_/A _22393_/X _21024_/X _22396_/X VGND VGND VPWR VPWR _22397_/X sky130_fd_sc_hd__a211o_4
X_12150_ _12104_/Y _12149_/X _12104_/Y _12149_/X VGND VGND VPWR VPWR _12157_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24136_ _24136_/CLK _18738_/X HRESETn VGND VGND VPWR VPWR _24136_/Q sky130_fd_sc_hd__dfrtp_4
X_21348_ _13533_/D _13789_/D _21344_/X _21559_/A _21347_/X VGND VGND VPWR VPWR _21348_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_123_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_118_0_HCLK clkbuf_7_59_0_HCLK/X VGND VGND VPWR VPWR _24561_/CLK sky130_fd_sc_hd__clkbuf_1
X_12081_ _12081_/A VGND VGND VPWR VPWR _12081_/Y sky130_fd_sc_hd__inv_2
X_24067_ _24069_/CLK _20526_/X HRESETn VGND VGND VPWR VPWR _20525_/A sky130_fd_sc_hd__dfrtp_4
X_21279_ _21859_/B VGND VGND VPWR VPWR _21280_/B sky130_fd_sc_hd__buf_2
XANTENNA__21149__B _21154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13530__A1 _13517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20760__A1_N _20743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23018_ _24589_/Q _22832_/B VGND VGND VPWR VPWR _23021_/B sky130_fd_sc_hd__or2_4
XFILLER_49_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15807__B1 _24830_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15840_ _14470_/A VGND VGND VPWR VPWR _15840_/X sky130_fd_sc_hd__buf_2
XFILLER_94_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17643__A _17525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16480__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15771_ _12562_/Y _15763_/X _14470_/X _15721_/A VGND VGND VPWR VPWR _24843_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15822__A3 _11809_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24496__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12983_ _12983_/A VGND VGND VPWR VPWR _13043_/A sky130_fd_sc_hd__inv_2
XANTENNA__12787__A _25357_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24969_ _24980_/CLK _15408_/X HRESETn VGND VGND VPWR VPWR _24969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21356__B2 _21549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17510_ _24302_/Q VGND VGND VPWR VPWR _17616_/A sky130_fd_sc_hd__inv_2
XFILLER_57_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20775__A1_N _20770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14722_ _14708_/X _14721_/X VGND VGND VPWR VPWR _14722_/X sky130_fd_sc_hd__or2_4
XFILLER_79_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11934_ _19615_/A VGND VGND VPWR VPWR _11934_/X sky130_fd_sc_hd__buf_2
X_18490_ _18496_/A _18490_/B VGND VGND VPWR VPWR _18503_/B sky130_fd_sc_hd__or2_4
XANTENNA__24425__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17441_ _14223_/B _21116_/A VGND VGND VPWR VPWR _17441_/Y sky130_fd_sc_hd__nor2_4
X_14653_ _17956_/A _14643_/Y VGND VGND VPWR VPWR _14653_/X sky130_fd_sc_hd__or2_4
X_11865_ HWDATA[0] VGND VGND VPWR VPWR _11865_/X sky130_fd_sc_hd__buf_2
X_13604_ _14645_/A _13610_/A VGND VGND VPWR VPWR _13605_/B sky130_fd_sc_hd__and2_4
XANTENNA__22708__B _21859_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17372_ _24333_/Q _17372_/B VGND VGND VPWR VPWR _17373_/C sky130_fd_sc_hd__or2_4
XANTENNA__14794__B1 _13598_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11796_ HWDATA[16] VGND VGND VPWR VPWR _11796_/X sky130_fd_sc_hd__buf_2
X_14584_ _14558_/X _14579_/B VGND VGND VPWR VPWR _14584_/X sky130_fd_sc_hd__or2_4
XFILLER_92_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19111_ _13263_/B VGND VGND VPWR VPWR _19111_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18193__B _18185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16323_ _16280_/X VGND VGND VPWR VPWR _16324_/A sky130_fd_sc_hd__buf_2
X_13535_ SSn_S2 _13534_/Y _13515_/X _13534_/Y VGND VGND VPWR VPWR _25291_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17732__B1 _21491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19042_ _23867_/Q VGND VGND VPWR VPWR _19042_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16254_ _16225_/A VGND VGND VPWR VPWR _16254_/X sky130_fd_sc_hd__buf_2
XANTENNA__15889__A3 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13466_ _15782_/B VGND VGND VPWR VPWR _15991_/B sky130_fd_sc_hd__buf_2
XFILLER_103_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15205_ _15069_/X _15171_/X _15070_/B VGND VGND VPWR VPWR _15205_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25284__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12417_ _12419_/B VGND VGND VPWR VPWR _12417_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12150__A1_N _12104_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16185_ _16373_/A _16459_/B VGND VGND VPWR VPWR _16192_/A sky130_fd_sc_hd__nor2_4
X_13397_ _13461_/A _13397_/B _13396_/X VGND VGND VPWR VPWR _13398_/C sky130_fd_sc_hd__or3_4
XANTENNA__16722__A _16722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_14_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__25213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15136_ _15135_/Y _24590_/Q _15135_/Y _24590_/Q VGND VGND VPWR VPWR _15141_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12348_ _12347_/Y _24819_/Q _12347_/Y _24819_/Q VGND VGND VPWR VPWR _12348_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_77_0_HCLK clkbuf_6_38_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_77_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11866__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12279_ _25430_/Q VGND VGND VPWR VPWR _12282_/C sky130_fd_sc_hd__inv_2
X_15067_ _15067_/A _15219_/B _15067_/C _15067_/D VGND VGND VPWR VPWR _15211_/A sky130_fd_sc_hd__or4_4
X_19944_ _19942_/Y _19943_/X _19629_/X _19943_/X VGND VGND VPWR VPWR _19944_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13784__C _13784_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14018_ _13977_/X _13980_/A _13984_/C _13983_/X VGND VGND VPWR VPWR _14018_/X sky130_fd_sc_hd__or4_4
X_19875_ _19875_/A VGND VGND VPWR VPWR _19875_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17553__A _17792_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18826_ _16537_/Y _24114_/Q _24539_/Q _18786_/C VGND VGND VPWR VPWR _18826_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18757_ _18757_/A _18757_/B VGND VGND VPWR VPWR _18758_/B sky130_fd_sc_hd__or2_4
XFILLER_97_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15969_ _15894_/A VGND VGND VPWR VPWR _15969_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17708_ _17708_/A VGND VGND VPWR VPWR _17708_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18688_ _18688_/A VGND VGND VPWR VPWR _18765_/A sky130_fd_sc_hd__inv_2
XFILLER_63_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17639_ _17564_/Y _17645_/B VGND VGND VPWR VPWR _17639_/X sky130_fd_sc_hd__or2_4
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12103__A1_N _12092_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20650_ _20650_/A _20650_/B VGND VGND VPWR VPWR _20650_/Y sky130_fd_sc_hd__nand2_4
X_19309_ _19309_/A VGND VGND VPWR VPWR _19309_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20858__B1 _20845_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20581_ _20580_/X VGND VGND VPWR VPWR _23941_/D sky130_fd_sc_hd__inv_2
XANTENNA__14417__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22320_ _23957_/Q VGND VGND VPWR VPWR _22320_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22251_ _22247_/A _22249_/X _22250_/X VGND VGND VPWR VPWR _22251_/X sky130_fd_sc_hd__and3_4
XANTENNA__12748__A1_N _25361_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21202_ _21201_/X VGND VGND VPWR VPWR _21202_/Y sky130_fd_sc_hd__inv_2
X_22182_ _21323_/A VGND VGND VPWR VPWR _22407_/B sky130_fd_sc_hd__buf_2
XFILLER_105_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21133_ _13517_/Y _21014_/A _13467_/X _21132_/Y VGND VGND VPWR VPWR _21133_/X sky130_fd_sc_hd__a211o_4
XANTENNA__11776__A _11776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19228__B1 _19136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21064_ _21064_/A VGND VGND VPWR VPWR _21064_/X sky130_fd_sc_hd__buf_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24936__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20015_ _20013_/Y _20014_/X _19992_/X _20014_/X VGND VGND VPWR VPWR _20015_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23184__B _21519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16462__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15804__A3 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24823_ _24821_/CLK _15818_/X HRESETn VGND VGND VPWR VPWR _24823_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12400__A _12385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24754_ _24759_/CLK _15961_/X HRESETn VGND VGND VPWR VPWR _22892_/A sky130_fd_sc_hd__dfrtp_4
X_21966_ _13775_/X _21965_/X VGND VGND VPWR VPWR _21966_/Y sky130_fd_sc_hd__nand2_4
XFILLER_104_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22809__A _22809_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23705_ _24926_/CLK _19503_/X VGND VGND VPWR VPWR _19502_/A sky130_fd_sc_hd__dfxtp_4
X_20917_ _20909_/X _20916_/Y _24488_/Q _20913_/X VGND VGND VPWR VPWR _20917_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _21622_/A _19918_/Y VGND VGND VPWR VPWR _21897_/X sky130_fd_sc_hd__or2_4
XPHY_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24685_ _24682_/CLK _24685_/D HRESETn VGND VGND VPWR VPWR _16122_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16807__A _16807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11650_/A VGND VGND VPWR VPWR _17445_/B sky130_fd_sc_hd__inv_2
XPHY_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _20846_/Y _20852_/B _20847_/X VGND VGND VPWR VPWR _20848_/X sky130_fd_sc_hd__o21a_4
XPHY_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23636_ _23635_/CLK _23636_/D VGND VGND VPWR VPWR _23636_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20329__A _20329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20849__B1 _20845_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20779_ _20779_/A VGND VGND VPWR VPWR _20779_/Y sky130_fd_sc_hd__inv_2
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23567_ _24309_/CLK _19903_/X VGND VGND VPWR VPWR _19901_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _13320_/A _23657_/Q VGND VGND VPWR VPWR _13320_/X sky130_fd_sc_hd__or2_4
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25306_ _25305_/CLK _25306_/D HRESETn VGND VGND VPWR VPWR _13488_/A sky130_fd_sc_hd__dfrtp_4
X_22518_ _22518_/A _22504_/Y _22511_/Y _22518_/D VGND VGND VPWR VPWR _22518_/X sky130_fd_sc_hd__or4_4
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23498_ _23498_/CLK _23498_/D VGND VGND VPWR VPWR _23498_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22544__A _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13251_ _13251_/A _13251_/B VGND VGND VPWR VPWR _13254_/B sky130_fd_sc_hd__or2_4
X_22449_ _22671_/A _22449_/B VGND VGND VPWR VPWR _22462_/A sky130_fd_sc_hd__nor2_4
X_25237_ _25192_/CLK _13870_/X HRESETn VGND VGND VPWR VPWR _22172_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_10_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16542__A _15709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12202_ _12202_/A VGND VGND VPWR VPWR _12282_/B sky130_fd_sc_hd__inv_2
X_13182_ _13186_/A _13182_/B VGND VGND VPWR VPWR _13182_/X sky130_fd_sc_hd__or2_4
X_25168_ _25305_/CLK _14298_/X HRESETn VGND VGND VPWR VPWR _13522_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11762__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12133_ _12125_/A _24096_/Q _12132_/Y VGND VGND VPWR VPWR _12134_/A sky130_fd_sc_hd__o21a_4
X_24119_ _24120_/CLK _18807_/X HRESETn VGND VGND VPWR VPWR _18601_/A sky130_fd_sc_hd__dfrtp_4
X_17990_ _17990_/A VGND VGND VPWR VPWR _18180_/A sky130_fd_sc_hd__buf_2
XANTENNA__23015__B2 _22827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25099_ _24077_/CLK _25099_/D HRESETn VGND VGND VPWR VPWR _20441_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12064_ _24914_/Q VGND VGND VPWR VPWR _16453_/A sky130_fd_sc_hd__buf_2
X_16941_ _16941_/A VGND VGND VPWR VPWR _16941_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24677__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19660_ _19660_/A VGND VGND VPWR VPWR _19660_/Y sky130_fd_sc_hd__inv_2
X_16872_ _16872_/A VGND VGND VPWR VPWR _16872_/X sky130_fd_sc_hd__buf_2
XANTENNA__23094__B _23075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24606__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18611_ _18610_/Y VGND VGND VPWR VPWR _18749_/A sky130_fd_sc_hd__buf_2
X_15823_ _15816_/X _15819_/X _15750_/X _24819_/Q _15817_/X VGND VGND VPWR VPWR _24819_/D
+ sky130_fd_sc_hd__a32o_4
X_19591_ _19590_/Y _19588_/X _19404_/X _19588_/X VGND VGND VPWR VPWR _19591_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17523__D _17522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18542_ _18461_/Y _18542_/B VGND VGND VPWR VPWR _18542_/Y sky130_fd_sc_hd__nand2_4
X_15754_ _15763_/A VGND VGND VPWR VPWR _15754_/X sky130_fd_sc_hd__buf_2
X_12966_ _25360_/Q _12966_/B VGND VGND VPWR VPWR _12967_/C sky130_fd_sc_hd__or2_4
XFILLER_79_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14705_ _14705_/A _14705_/B VGND VGND VPWR VPWR _14705_/X sky130_fd_sc_hd__or2_4
X_11917_ _11876_/X _11902_/B VGND VGND VPWR VPWR _11917_/Y sky130_fd_sc_hd__nor2_4
X_18473_ _24149_/Q VGND VGND VPWR VPWR _18475_/B sky130_fd_sc_hd__inv_2
X_15685_ _15685_/A VGND VGND VPWR VPWR _15685_/X sky130_fd_sc_hd__buf_2
X_12897_ _12881_/A _12887_/X _12897_/C VGND VGND VPWR VPWR _12897_/X sky130_fd_sc_hd__and3_4
XANTENNA__16717__A _14470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17424_ _16528_/A VGND VGND VPWR VPWR _17424_/X sky130_fd_sc_hd__buf_2
X_14636_ _18079_/A VGND VGND VPWR VPWR _18059_/A sky130_fd_sc_hd__buf_2
XANTENNA__22829__A1 _23126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11848_ _11750_/A VGND VGND VPWR VPWR _11848_/X sky130_fd_sc_hd__buf_2
XANTENNA__25465__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17355_ _17350_/A _17350_/B _17349_/X VGND VGND VPWR VPWR _17355_/X sky130_fd_sc_hd__or3_4
X_14567_ _13576_/Y _14567_/B VGND VGND VPWR VPWR _14592_/B sky130_fd_sc_hd__or2_4
X_11779_ _11776_/Y _11777_/X _11778_/X _11777_/X VGND VGND VPWR VPWR _25528_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16306_ HWDATA[23] VGND VGND VPWR VPWR _16306_/X sky130_fd_sc_hd__buf_2
XFILLER_105_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13518_ _13517_/Y _13512_/X _13472_/X _13512_/X VGND VGND VPWR VPWR _25294_/D sky130_fd_sc_hd__a2bb2o_4
X_17286_ _17266_/A _17286_/B _17285_/X VGND VGND VPWR VPWR _17286_/X sky130_fd_sc_hd__and3_4
X_14498_ _14497_/X VGND VGND VPWR VPWR _14498_/Y sky130_fd_sc_hd__inv_2
X_19025_ _23873_/Q VGND VGND VPWR VPWR _19025_/Y sky130_fd_sc_hd__inv_2
X_16237_ _22619_/A VGND VGND VPWR VPWR _16237_/Y sky130_fd_sc_hd__inv_2
X_13449_ _13417_/A _19702_/A VGND VGND VPWR VPWR _13450_/C sky130_fd_sc_hd__or2_4
XANTENNA__23254__A1 _21409_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16168_ _16173_/A _14770_/B VGND VGND VPWR VPWR _16169_/A sky130_fd_sc_hd__or2_4
XANTENNA__13795__B _16725_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15119_ _24981_/Q _24585_/Q _15367_/A _15118_/Y VGND VGND VPWR VPWR _15120_/D sky130_fd_sc_hd__o22a_4
XANTENNA__23006__A1 _24524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16099_ _16098_/Y _16094_/X _15944_/X _16094_/X VGND VGND VPWR VPWR _16099_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19927_ _23557_/Q VGND VGND VPWR VPWR _19927_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_101_0_HCLK clkbuf_7_50_0_HCLK/X VGND VGND VPWR VPWR _24151_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_130_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_164_0_HCLK clkbuf_7_82_0_HCLK/X VGND VGND VPWR VPWR _23598_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24347__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_7_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19858_ _19858_/A VGND VGND VPWR VPWR _19858_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18433__B2 _24168_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16444__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18809_ _18809_/A _18809_/B VGND VGND VPWR VPWR _18810_/C sky130_fd_sc_hd__or2_4
X_19789_ _19789_/A VGND VGND VPWR VPWR _21748_/B sky130_fd_sc_hd__inv_2
X_21820_ _13784_/D _21819_/X VGND VGND VPWR VPWR _21820_/X sky130_fd_sc_hd__or2_4
XFILLER_83_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21751_ _21747_/X _21750_/X _14712_/X VGND VGND VPWR VPWR _21751_/X sky130_fd_sc_hd__o21a_4
XFILLER_3_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21533__A _21418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21740__A1 _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20702_ _20702_/A VGND VGND VPWR VPWR _20702_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15531__A _11726_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21682_ _21661_/X _21681_/X _21493_/X VGND VGND VPWR VPWR _21682_/Y sky130_fd_sc_hd__a21oi_4
X_24470_ _24035_/CLK _24470_/D HRESETn VGND VGND VPWR VPWR _24470_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23982__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20633_ _20633_/A _17392_/X VGND VGND VPWR VPWR _20635_/B sky130_fd_sc_hd__nand2_4
XFILLER_75_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23421_ _23398_/CLK _23421_/D VGND VGND VPWR VPWR _23421_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22296__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25135__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23352_ VGND VGND VPWR VPWR _23352_/HI sda_o_S4 sky130_fd_sc_hd__conb_1
X_20564_ _14430_/Y _20556_/X _20547_/X _20563_/X VGND VGND VPWR VPWR _20565_/A sky130_fd_sc_hd__a211o_4
XFILLER_137_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22303_ _14373_/Y _14192_/X _14474_/Y _21139_/B VGND VGND VPWR VPWR _22304_/A sky130_fd_sc_hd__o22a_4
X_23283_ _17235_/Y _22475_/X _12830_/A _22435_/X VGND VGND VPWR VPWR _23283_/X sky130_fd_sc_hd__a2bb2o_4
X_20495_ _14063_/X _20439_/X VGND VGND VPWR VPWR _20495_/X sky130_fd_sc_hd__and2_4
XANTENNA__12890__A _12749_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22234_ _22229_/A _22234_/B VGND VGND VPWR VPWR _22234_/X sky130_fd_sc_hd__or2_4
X_25022_ _25020_/CLK _15188_/X HRESETn VGND VGND VPWR VPWR _25022_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16081__B _15674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11744__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22165_ _22158_/Y _22160_/Y _22163_/Y _22164_/X VGND VGND VPWR VPWR _22165_/X sky130_fd_sc_hd__or4_4
XFILLER_65_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_60_0_HCLK clkbuf_6_30_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21116_ _21116_/A VGND VGND VPWR VPWR _21116_/Y sky130_fd_sc_hd__inv_2
X_22096_ _22095_/X VGND VGND VPWR VPWR _22101_/B sky130_fd_sc_hd__inv_2
XANTENNA__24770__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21047_ _21306_/A VGND VGND VPWR VPWR _21048_/B sky130_fd_sc_hd__buf_2
XANTENNA__15706__A _21154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24088__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16435__B1 _16064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24017__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16986__A1 _24705_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12820_ _23213_/A VGND VGND VPWR VPWR _12820_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13226__A _13310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24806_ _24806_/CLK _15844_/X HRESETn VGND VGND VPWR VPWR _21006_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_28_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22998_ _22998_/A VGND VGND VPWR VPWR _22998_/X sky130_fd_sc_hd__buf_2
XANTENNA__21825__A2_N _21306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12751_ _12743_/X _12745_/X _12751_/C _12750_/X VGND VGND VPWR VPWR _12791_/A sky130_fd_sc_hd__or4_4
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24737_ _24792_/CLK _15987_/X HRESETn VGND VGND VPWR VPWR _21526_/A sky130_fd_sc_hd__dfrtp_4
X_21949_ _21160_/X VGND VGND VPWR VPWR _21950_/A sky130_fd_sc_hd__buf_2
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16537__A _24535_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11961_/A _11967_/D _11702_/C VGND VGND VPWR VPWR _11970_/D sky130_fd_sc_hd__and3_4
XFILLER_76_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15470_/A VGND VGND VPWR VPWR _15470_/Y sky130_fd_sc_hd__inv_2
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12686_/A _12682_/B _12682_/C VGND VGND VPWR VPWR _25406_/D sky130_fd_sc_hd__and3_4
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24668_ _24606_/CLK _24668_/D HRESETn VGND VGND VPWR VPWR _21051_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _25129_/Q VGND VGND VPWR VPWR _14421_/Y sky130_fd_sc_hd__inv_2
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ _23635_/CLK _23619_/D VGND VGND VPWR VPWR _13251_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24599_ _24889_/CLK _16367_/X HRESETn VGND VGND VPWR VPWR _24599_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17140_ _17038_/A _17134_/B VGND VGND VPWR VPWR _17141_/C sky130_fd_sc_hd__nand2_4
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14352_ _14339_/Y _14336_/C _14325_/X _14351_/X VGND VGND VPWR VPWR _14353_/A sky130_fd_sc_hd__a211o_4
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _13303_/A _13303_/B VGND VGND VPWR VPWR _13303_/X sky130_fd_sc_hd__or2_4
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17071_ _24387_/Q _17071_/B VGND VGND VPWR VPWR _17073_/B sky130_fd_sc_hd__or2_4
X_14283_ _20467_/A _14281_/X _20467_/A _14282_/X VGND VGND VPWR VPWR _14283_/X sky130_fd_sc_hd__o22a_4
XFILLER_13_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16022_ _16002_/X VGND VGND VPWR VPWR _16022_/X sky130_fd_sc_hd__buf_2
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13234_ _13234_/A VGND VGND VPWR VPWR _13455_/A sky130_fd_sc_hd__buf_2
XFILLER_13_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24858__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13165_ _13180_/A VGND VGND VPWR VPWR _13190_/A sky130_fd_sc_hd__buf_2
XANTENNA__19860__B1 _19794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12305__A _12305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25126__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16674__B1 _16405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12116_ _12116_/A VGND VGND VPWR VPWR _12116_/Y sky130_fd_sc_hd__inv_2
X_13096_ _13096_/A _13084_/B VGND VGND VPWR VPWR _13096_/Y sky130_fd_sc_hd__nand2_4
X_17973_ _17996_/A VGND VGND VPWR VPWR _17973_/X sky130_fd_sc_hd__buf_2
XANTENNA__21618__A _21618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12047_ _16371_/A VGND VGND VPWR VPWR _16183_/A sky130_fd_sc_hd__buf_2
X_16924_ _17826_/A VGND VGND VPWR VPWR _17758_/B sky130_fd_sc_hd__inv_2
X_19712_ _19706_/Y VGND VGND VPWR VPWR _19712_/X sky130_fd_sc_hd__buf_2
XANTENNA__18415__A1 _23242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18415__B2 _18481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24440__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18432__A1_N _16234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_237_0_HCLK clkbuf_8_237_0_HCLK/A VGND VGND VPWR VPWR _24836_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_93_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16855_ _16855_/A VGND VGND VPWR VPWR _16855_/Y sky130_fd_sc_hd__inv_2
X_19643_ _19641_/Y _19639_/X _19642_/X _19639_/X VGND VGND VPWR VPWR _23659_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15806_ _12321_/Y _15802_/X _11767_/X _15802_/X VGND VGND VPWR VPWR _15806_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21970__B2 _21636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19574_ _19574_/A VGND VGND VPWR VPWR _19574_/X sky130_fd_sc_hd__buf_2
XANTENNA__11849__A1_N _11844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16786_ HWDATA[3] VGND VGND VPWR VPWR _16786_/X sky130_fd_sc_hd__buf_2
X_13998_ _13990_/B VGND VGND VPWR VPWR _13998_/X sky130_fd_sc_hd__buf_2
XFILLER_46_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22449__A _22671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18525_ _18525_/A VGND VGND VPWR VPWR _18525_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15737_ _12555_/Y _15735_/X _11788_/X _15735_/X VGND VGND VPWR VPWR _24860_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18447__A1_N _23232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12949_ _12955_/A _12944_/B _12944_/D VGND VGND VPWR VPWR _12949_/X sky130_fd_sc_hd__or3_4
XANTENNA__21722__B2 _16723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15351__A _15336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18456_ _18456_/A _18503_/A VGND VGND VPWR VPWR _18456_/X sky130_fd_sc_hd__or2_4
X_15668_ _15668_/A VGND VGND VPWR VPWR _15668_/X sky130_fd_sc_hd__buf_2
X_17407_ _17387_/X _17401_/X _23986_/Q _20992_/B _17404_/X VGND VGND VPWR VPWR _24325_/D
+ sky130_fd_sc_hd__a32o_4
X_14619_ _14619_/A VGND VGND VPWR VPWR _14620_/A sky130_fd_sc_hd__inv_2
X_18387_ _18386_/Y _18384_/X _24178_/Q _18384_/X VGND VGND VPWR VPWR _18387_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19679__B1 _19462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19758__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15599_ _15599_/A VGND VGND VPWR VPWR _15599_/Y sky130_fd_sc_hd__inv_2
X_17338_ _17337_/X VGND VGND VPWR VPWR _17338_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22184__A _21859_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17269_ _17194_/Y _17261_/B _17269_/C VGND VGND VPWR VPWR _17269_/X sky130_fd_sc_hd__or3_4
XFILLER_119_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19008_ _19007_/Y _19005_/X _18940_/X _19005_/X VGND VGND VPWR VPWR _23878_/D sky130_fd_sc_hd__a2bb2o_4
X_20280_ _23426_/Q VGND VGND VPWR VPWR _22250_/B sky130_fd_sc_hd__inv_2
XANTENNA__24599__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24528__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22631__B _23035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_47_0_HCLK clkbuf_6_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16665__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22738__B1 _24857_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24181__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19603__B1 _19553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14430__A _25125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23970_ _24942_/CLK _23970_/D HRESETn VGND VGND VPWR VPWR _17388_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_69_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16417__B1 _16228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22921_ _16216_/A _22796_/B VGND VGND VPWR VPWR _22926_/B sky130_fd_sc_hd__or2_4
XFILLER_96_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20764__A2 _20676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22852_ _22814_/X _22818_/X _22852_/C _22851_/X VGND VGND VPWR VPWR HRDATA[17] sky130_fd_sc_hd__or4_4
XFILLER_43_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_21803_ _21477_/A _21803_/B VGND VGND VPWR VPWR _21803_/X sky130_fd_sc_hd__or2_4
XANTENNA__25387__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22783_ _22783_/A VGND VGND VPWR VPWR _22783_/X sky130_fd_sc_hd__buf_2
XANTENNA__25316__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24522_ _24555_/CLK _24522_/D HRESETn VGND VGND VPWR VPWR _24522_/Q sky130_fd_sc_hd__dfrtp_4
X_21734_ _16533_/Y _22695_/C VGND VGND VPWR VPWR _21734_/X sky130_fd_sc_hd__and2_4
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24453_ _25024_/CLK _24453_/D HRESETn VGND VGND VPWR VPWR _24453_/Q sky130_fd_sc_hd__dfrtp_4
X_21665_ _21670_/A _20310_/Y VGND VGND VPWR VPWR _21665_/X sky130_fd_sc_hd__or2_4
XFILLER_36_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23404_ _24208_/CLK _23404_/D VGND VGND VPWR VPWR _20335_/A sky130_fd_sc_hd__dfxtp_4
X_20616_ _15470_/Y _20605_/X _20662_/A _20615_/X VGND VGND VPWR VPWR _20617_/A sky130_fd_sc_hd__a211o_4
X_21596_ _21596_/A _19835_/Y VGND VGND VPWR VPWR _21599_/B sky130_fd_sc_hd__or2_4
X_24384_ _24368_/CLK _17083_/X HRESETn VGND VGND VPWR VPWR _24384_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20547_ _20546_/X VGND VGND VPWR VPWR _20547_/X sky130_fd_sc_hd__buf_2
X_23335_ _23334_/X VGND VGND VPWR VPWR _23335_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20478_ _24070_/Q _20502_/A VGND VGND VPWR VPWR _20479_/C sky130_fd_sc_hd__and2_4
XANTENNA__24951__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23266_ _23265_/X VGND VGND VPWR VPWR _23266_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22977__B1 _11776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25005_ _25001_/CLK _15258_/Y HRESETn VGND VGND VPWR VPWR _25005_/Q sky130_fd_sc_hd__dfrtp_4
X_22217_ _21601_/A _22215_/X _22216_/X VGND VGND VPWR VPWR _22218_/C sky130_fd_sc_hd__and3_4
XFILLER_69_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19842__B1 _19841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24269__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23197_ _23124_/A _23197_/B VGND VGND VPWR VPWR _23197_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__16656__B1 _16297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22148_ _22134_/X _22148_/B VGND VGND VPWR VPWR _22148_/X sky130_fd_sc_hd__and2_4
XANTENNA__21438__A _21009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14970_ _15071_/A _24427_/Q _25015_/Q _14969_/Y VGND VGND VPWR VPWR _14970_/X sky130_fd_sc_hd__a2bb2o_4
X_22079_ _22070_/X _19851_/Y _22078_/X VGND VGND VPWR VPWR _22079_/X sky130_fd_sc_hd__o21a_4
XFILLER_134_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13921_ _13945_/A VGND VGND VPWR VPWR _13921_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16640_ _16640_/A _16640_/B VGND VGND VPWR VPWR _16643_/A sky130_fd_sc_hd__or2_4
XFILLER_74_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13852_ _23989_/Q VGND VGND VPWR VPWR _13852_/X sky130_fd_sc_hd__buf_2
XFILLER_16_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_67_0_HCLK clkbuf_8_67_0_HCLK/A VGND VGND VPWR VPWR _25137_/CLK sky130_fd_sc_hd__clkbuf_1
X_12803_ _12924_/A _22708_/A _12924_/A _22708_/A VGND VGND VPWR VPWR _12803_/X sky130_fd_sc_hd__a2bb2o_4
X_16571_ _16569_/Y _16570_/X _16401_/X _16570_/X VGND VGND VPWR VPWR _16571_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13783_ _13782_/X VGND VGND VPWR VPWR _13784_/D sky130_fd_sc_hd__buf_2
X_18310_ _21658_/A _18300_/A _18303_/X VGND VGND VPWR VPWR _24199_/D sky130_fd_sc_hd__a21oi_4
X_15522_ _15521_/Y _15517_/X HADDR[10] _15517_/X VGND VGND VPWR VPWR _24922_/D sky130_fd_sc_hd__a2bb2o_4
X_12734_ _12731_/B _12734_/B _12721_/X VGND VGND VPWR VPWR _12734_/X sky130_fd_sc_hd__and3_4
X_19290_ _13240_/B VGND VGND VPWR VPWR _19290_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18241_ _18235_/X _18237_/X _11812_/X _24225_/Q _18238_/X VGND VGND VPWR VPWR _18241_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_37_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15453_ _13905_/C _15449_/X _15446_/X _13901_/X _15452_/X VGND VGND VPWR VPWR _15453_/X
+ sky130_fd_sc_hd__a32o_4
X_12665_ _12665_/A _12618_/X VGND VGND VPWR VPWR _12674_/B sky130_fd_sc_hd__or2_4
XFILLER_54_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _20592_/A _14384_/A _14403_/X _14384_/A VGND VGND VPWR VPWR _25133_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21468__B1 _18299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18172_ _18204_/A _18172_/B VGND VGND VPWR VPWR _18172_/X sky130_fd_sc_hd__or2_4
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15384_ _15384_/A _15384_/B _15384_/C VGND VGND VPWR VPWR _24976_/D sky130_fd_sc_hd__and3_4
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _12596_/A VGND VGND VPWR VPWR _12731_/A sky130_fd_sc_hd__buf_2
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11956__B1 _11955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17123_ _17036_/Y _17120_/X VGND VGND VPWR VPWR _17123_/X sky130_fd_sc_hd__or2_4
X_14335_ _18370_/B _14333_/X VGND VGND VPWR VPWR _14336_/C sky130_fd_sc_hd__or2_4
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17054_ _17064_/A _17052_/X _17054_/C VGND VGND VPWR VPWR _17054_/X sky130_fd_sc_hd__and3_4
XFILLER_7_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14266_ _14266_/A VGND VGND VPWR VPWR _14266_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24692__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16005_ _24731_/Q VGND VGND VPWR VPWR _16005_/Y sky130_fd_sc_hd__inv_2
X_13217_ _13162_/A VGND VGND VPWR VPWR _13314_/A sky130_fd_sc_hd__buf_2
XANTENNA__24621__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14197_ _20657_/A VGND VGND VPWR VPWR _14807_/A sky130_fd_sc_hd__inv_2
XFILLER_48_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16647__B1 _16285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13148_ _13251_/A VGND VGND VPWR VPWR _13186_/A sky130_fd_sc_hd__buf_2
XFILLER_48_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13079_ _12311_/Y _13043_/A VGND VGND VPWR VPWR _13113_/A sky130_fd_sc_hd__or2_4
X_17956_ _17956_/A _23892_/Q VGND VGND VPWR VPWR _17957_/C sky130_fd_sc_hd__or2_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16907_ _24253_/Q VGND VGND VPWR VPWR _17846_/A sky130_fd_sc_hd__inv_2
XFILLER_66_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17887_ _24244_/Q VGND VGND VPWR VPWR _17887_/Y sky130_fd_sc_hd__inv_2
X_19626_ _21811_/B _19619_/X _19625_/X _19619_/X VGND VGND VPWR VPWR _19626_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16838_ _16836_/Y _16837_/X _15752_/X _16837_/X VGND VGND VPWR VPWR _24412_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23145__B1 _24868_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21083__A _21024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25480__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16769_ _24444_/Q VGND VGND VPWR VPWR _16769_/Y sky130_fd_sc_hd__inv_2
X_19557_ _23685_/Q VGND VGND VPWR VPWR _19557_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22499__A2 _22444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18508_ _16448_/A _18478_/B _18442_/Y _18466_/X VGND VGND VPWR VPWR _18508_/X sky130_fd_sc_hd__or4_4
XFILLER_34_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19488_ _19885_/A VGND VGND VPWR VPWR _19488_/X sky130_fd_sc_hd__buf_2
XFILLER_62_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18439_ _16258_/Y _24149_/Q _23232_/A _18456_/A VGND VGND VPWR VPWR _18439_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22626__B _22626_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21450_ _21478_/A VGND VGND VPWR VPWR _21648_/A sky130_fd_sc_hd__buf_2
X_20401_ _20397_/Y _20400_/X _18247_/X _20400_/X VGND VGND VPWR VPWR _20401_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_4_10_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_10_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_21381_ _21381_/A _21381_/B VGND VGND VPWR VPWR _21381_/X sky130_fd_sc_hd__or2_4
XANTENNA__24709__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20332_ _20331_/Y _20327_/X _20072_/X _20327_/X VGND VGND VPWR VPWR _23406_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23120_ _23120_/A _22914_/B VGND VGND VPWR VPWR _23120_/X sky130_fd_sc_hd__and2_4
X_23051_ _16662_/Y _22914_/B VGND VGND VPWR VPWR _23051_/X sky130_fd_sc_hd__and2_4
X_20263_ _23432_/Q VGND VGND VPWR VPWR _21769_/B sky130_fd_sc_hd__inv_2
XANTENNA__23223__A2_N _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24362__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22423__A2 _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16640__A _16640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22002_ _22247_/A VGND VGND VPWR VPWR _22025_/A sky130_fd_sc_hd__buf_2
XFILLER_88_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20194_ _22216_/B _20191_/X _19780_/A _20191_/X VGND VGND VPWR VPWR _20194_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23176__C _23169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11784__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12124__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23953_ _25219_/CLK _20598_/X HRESETn VGND VGND VPWR VPWR _23953_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_220_0_HCLK clkbuf_8_221_0_HCLK/A VGND VGND VPWR VPWR _25002_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_29_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22904_ _22769_/X _22901_/Y _22863_/X _22903_/X VGND VGND VPWR VPWR _22904_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23884_ _23884_/CLK _23884_/D VGND VGND VPWR VPWR _23884_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23136__B1 _22997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22089__A _22089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16810__B1 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18286__B _17702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22835_ _22835_/A VGND VGND VPWR VPWR _23019_/C sky130_fd_sc_hd__buf_2
XANTENNA__21698__B1 _24810_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25150__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22766_ _21418_/X VGND VGND VPWR VPWR _22766_/X sky130_fd_sc_hd__buf_2
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24505_ _24545_/CLK _16617_/X HRESETn VGND VGND VPWR VPWR _16616_/A sky130_fd_sc_hd__dfrtp_4
X_21717_ _21716_/Y _21143_/X _15473_/Y _21352_/X VGND VGND VPWR VPWR _21718_/A sky130_fd_sc_hd__o22a_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15916__A2 _13588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25485_ _25485_/CLK _25485_/D HRESETn VGND VGND VPWR VPWR _11654_/C sky130_fd_sc_hd__dfrtp_4
X_22697_ _23085_/A _22694_/X _22696_/X VGND VGND VPWR VPWR _22711_/A sky130_fd_sc_hd__and3_4
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17533__A1_N _11807_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _12440_/C _12432_/B _12402_/X _12448_/B VGND VGND VPWR VPWR _12451_/A sky130_fd_sc_hd__a211o_4
X_24436_ _24435_/CLK _16788_/X HRESETn VGND VGND VPWR VPWR _16785_/A sky130_fd_sc_hd__dfrtp_4
X_21648_ _21648_/A _20289_/Y VGND VGND VPWR VPWR _21649_/C sky130_fd_sc_hd__or2_4
XANTENNA__11959__A _11958_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ _12351_/X _12381_/B _12381_/C _12380_/X VGND VGND VPWR VPWR _12382_/B sky130_fd_sc_hd__or4_4
X_24367_ _24368_/CLK _17145_/X HRESETn VGND VGND VPWR VPWR _24367_/Q sky130_fd_sc_hd__dfrtp_4
X_21579_ _21281_/X VGND VGND VPWR VPWR _21580_/A sky130_fd_sc_hd__buf_2
XANTENNA__18866__B2 _18865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14120_ _14106_/C _14120_/B VGND VGND VPWR VPWR _14120_/Y sky130_fd_sc_hd__nor2_4
X_23318_ _23318_/A _16795_/A VGND VGND VPWR VPWR _23318_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24311__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24298_ _25526_/CLK _17633_/Y HRESETn VGND VGND VPWR VPWR _24298_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13596__D _13777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17548__A1_N _11753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14051_ _14070_/A _14543_/C _14038_/Y _14050_/X VGND VGND VPWR VPWR _14051_/X sky130_fd_sc_hd__or4_4
XFILLER_101_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18618__A1 _24520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23249_ _22646_/A _23246_/X _23248_/X VGND VGND VPWR VPWR _23249_/X sky130_fd_sc_hd__and3_4
X_13002_ _12374_/Y _13002_/B _13001_/X VGND VGND VPWR VPWR _13005_/B sky130_fd_sc_hd__or3_4
XFILLER_136_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24032__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20072__A _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_30_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_30_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17810_ _17758_/X _17818_/D VGND VGND VPWR VPWR _17810_/X sky130_fd_sc_hd__or2_4
XFILLER_0_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18790_ _18680_/A _18788_/A VGND VGND VPWR VPWR _18791_/C sky130_fd_sc_hd__or2_4
XANTENNA__12115__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17741_ _24268_/Q VGND VGND VPWR VPWR _17741_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14953_ _15068_/A VGND VGND VPWR VPWR _15209_/A sky130_fd_sc_hd__buf_2
XFILLER_48_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13904_ _24950_/Q VGND VGND VPWR VPWR _13904_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25238__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17672_ _17499_/Y _17672_/B VGND VGND VPWR VPWR _17672_/Y sky130_fd_sc_hd__nand2_4
X_14884_ pwm_S6 VGND VGND VPWR VPWR _14884_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16623_ _16622_/Y _16545_/A _16366_/X _16545_/A VGND VGND VPWR VPWR _16623_/X sky130_fd_sc_hd__a2bb2o_4
X_19411_ _19410_/Y _19408_/X _19364_/X _19408_/X VGND VGND VPWR VPWR _23737_/D sky130_fd_sc_hd__a2bb2o_4
X_13835_ _13835_/A VGND VGND VPWR VPWR _13835_/X sky130_fd_sc_hd__buf_2
XFILLER_112_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13414__A _13162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16554_ _16553_/Y _16551_/X _16384_/X _16551_/X VGND VGND VPWR VPWR _24530_/D sky130_fd_sc_hd__a2bb2o_4
X_19342_ _19341_/Y _19339_/X _19206_/X _19339_/X VGND VGND VPWR VPWR _23761_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13766_ _13752_/A VGND VGND VPWR VPWR _20043_/D sky130_fd_sc_hd__buf_2
XFILLER_56_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21153__A2 _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22350__A1 _17706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15505_ _15503_/Y _15499_/X HADDR[17] _15504_/X VGND VGND VPWR VPWR _24929_/D sky130_fd_sc_hd__a2bb2o_4
X_12717_ _12698_/A _12708_/B _12716_/Y VGND VGND VPWR VPWR _12717_/X sky130_fd_sc_hd__and3_4
X_19273_ _19273_/A VGND VGND VPWR VPWR _21886_/B sky130_fd_sc_hd__inv_2
X_16485_ _16485_/A VGND VGND VPWR VPWR _16485_/Y sky130_fd_sc_hd__inv_2
X_13697_ _13676_/Y _13680_/X _13693_/X _13676_/A _13696_/Y VGND VGND VPWR VPWR _13697_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16725__A _16725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18224_ _18224_/A _18224_/B _18223_/X VGND VGND VPWR VPWR _18224_/X sky130_fd_sc_hd__or3_4
X_15436_ _13952_/A _15432_/X _15435_/X VGND VGND VPWR VPWR _15436_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21350__B _21350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12648_ _12648_/A _12644_/B _12647_/X VGND VGND VPWR VPWR _12648_/X sky130_fd_sc_hd__or3_4
XANTENNA__24873__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18155_ _18187_/A _19166_/A VGND VGND VPWR VPWR _18156_/C sky130_fd_sc_hd__or2_4
X_15367_ _15367_/A _15370_/B VGND VGND VPWR VPWR _15368_/C sky130_fd_sc_hd__nand2_4
XANTENNA__24802__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12579_ _25410_/Q VGND VGND VPWR VPWR _12620_/B sky130_fd_sc_hd__inv_2
XFILLER_102_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18940__A _14470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17106_ _17034_/B _17105_/X VGND VGND VPWR VPWR _17110_/B sky130_fd_sc_hd__or2_4
XFILLER_116_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14318_ _14305_/Y _14317_/X _25307_/Q _14311_/X VGND VGND VPWR VPWR _25161_/D sky130_fd_sc_hd__o22a_4
X_18086_ _18185_/A _18086_/B _18086_/C VGND VGND VPWR VPWR _18097_/B sky130_fd_sc_hd__or3_4
XFILLER_8_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15298_ _15356_/A _15298_/B _15298_/C VGND VGND VPWR VPWR _15336_/D sky130_fd_sc_hd__or3_4
Xclkbuf_7_112_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_225_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17037_ _24372_/Q VGND VGND VPWR VPWR _17120_/A sky130_fd_sc_hd__inv_2
X_14249_ _14249_/A _13931_/Y VGND VGND VPWR VPWR _15428_/A sky130_fd_sc_hd__or2_4
XANTENNA__17556__A _24308_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19806__B1 _19755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22181__B _21220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21078__A _15852_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19771__A _15845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18988_ _18987_/X VGND VGND VPWR VPWR _18988_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17939_ _14648_/X _17939_/B _17939_/C VGND VGND VPWR VPWR _17939_/X sky130_fd_sc_hd__and3_4
XFILLER_117_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20950_ _20812_/A _24060_/Q _13667_/X _23317_/A _20864_/X VGND VGND VPWR VPWR _24060_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_96_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19609_ _18275_/X _20338_/B _20276_/C VGND VGND VPWR VPWR _19609_/X sky130_fd_sc_hd__or3_4
X_20881_ _20860_/X _20880_/X _24480_/Q _20865_/X VGND VGND VPWR VPWR _20881_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_50_0_HCLK clkbuf_8_51_0_HCLK/A VGND VGND VPWR VPWR _25070_/CLK sky130_fd_sc_hd__clkbuf_1
X_22620_ _16508_/A _22422_/X _22527_/X VGND VGND VPWR VPWR _22620_/X sky130_fd_sc_hd__o21a_4
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21144__A2 _14192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21541__A _21333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22551_ _21111_/X VGND VGND VPWR VPWR _22551_/X sky130_fd_sc_hd__buf_2
XANTENNA__21695__A3 _21514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21502_ _21502_/A VGND VGND VPWR VPWR _21502_/X sky130_fd_sc_hd__buf_2
XFILLER_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25270_ _24214_/CLK _25270_/D HRESETn VGND VGND VPWR VPWR _25270_/Q sky130_fd_sc_hd__dfrtp_4
X_22482_ _22482_/A VGND VGND VPWR VPWR _22482_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24221_ _24715_/CLK _24221_/D HRESETn VGND VGND VPWR VPWR _24221_/Q sky130_fd_sc_hd__dfrtp_4
X_21433_ _21433_/A _22590_/B VGND VGND VPWR VPWR _21433_/X sky130_fd_sc_hd__or2_4
XFILLER_108_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24543__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21364_ _21996_/A _19536_/Y _21364_/C VGND VGND VPWR VPWR _21499_/B sky130_fd_sc_hd__or3_4
X_24152_ _24643_/CLK _24152_/D HRESETn VGND VGND VPWR VPWR _24152_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17520__A1 _25509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20315_ _20315_/A VGND VGND VPWR VPWR _21164_/B sky130_fd_sc_hd__inv_2
X_23103_ _23034_/X _23101_/X _22968_/X _24867_/Q _23102_/X VGND VGND VPWR VPWR _23104_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_107_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21295_ _22138_/A VGND VGND VPWR VPWR _21295_/X sky130_fd_sc_hd__buf_2
X_24083_ _23847_/CLK _20951_/X HRESETn VGND VGND VPWR VPWR RsTx_S1 sky130_fd_sc_hd__dfstp_4
XANTENNA__16370__A _16722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20246_ _20244_/Y _20245_/X _20072_/X _20245_/X VGND VGND VPWR VPWR _23439_/D sky130_fd_sc_hd__a2bb2o_4
X_23034_ _23034_/A VGND VGND VPWR VPWR _23034_/X sky130_fd_sc_hd__buf_2
XFILLER_27_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_17_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20177_ _23465_/Q VGND VGND VPWR VPWR _20177_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18831__A1_N _16533_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13845__B1 _13803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24985_ _24984_/CLK _24985_/D HRESETn VGND VGND VPWR VPWR _24985_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15714__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25331__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11950_ _19995_/A VGND VGND VPWR VPWR _19632_/A sky130_fd_sc_hd__buf_2
X_23936_ _24364_/CLK _23936_/D HRESETn VGND VGND VPWR VPWR _18874_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15598__B1 _11796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11881_ _11880_/Y VGND VGND VPWR VPWR _13678_/B sky130_fd_sc_hd__buf_2
X_23867_ _25485_/CLK _19043_/X VGND VGND VPWR VPWR _23867_/Q sky130_fd_sc_hd__dfxtp_4
X_13620_ _13619_/X VGND VGND VPWR VPWR _14661_/A sky130_fd_sc_hd__inv_2
X_22818_ _22270_/X _22815_/X _22817_/X VGND VGND VPWR VPWR _22818_/X sky130_fd_sc_hd__and3_4
X_23798_ _23798_/CLK _19238_/X VGND VGND VPWR VPWR _13404_/B sky130_fd_sc_hd__dfxtp_4
X_13551_ _13551_/A VGND VGND VPWR VPWR _13551_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25537_ _24267_/CLK _11747_/X HRESETn VGND VGND VPWR VPWR _25537_/Q sky130_fd_sc_hd__dfrtp_4
X_22749_ _22827_/A _22747_/X _22103_/X _22748_/X VGND VGND VPWR VPWR _22750_/B sky130_fd_sc_hd__o22a_4
XFILLER_125_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16545__A _16545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12502_ _12499_/A _12499_/B VGND VGND VPWR VPWR _12502_/Y sky130_fd_sc_hd__nand2_4
X_16270_ _11865_/X VGND VGND VPWR VPWR _16270_/X sky130_fd_sc_hd__buf_2
XFILLER_73_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13482_ _13476_/Y VGND VGND VPWR VPWR _13482_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25468_ _24097_/CLK _25468_/D HRESETn VGND VGND VPWR VPWR _25468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15221_ _14926_/X _15219_/X _15220_/Y VGND VGND VPWR VPWR _25014_/D sky130_fd_sc_hd__o21a_4
X_12433_ _12433_/A _12433_/B VGND VGND VPWR VPWR _12433_/X sky130_fd_sc_hd__or2_4
X_24419_ _24431_/CLK _24419_/D HRESETn VGND VGND VPWR VPWR _14913_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15770__B1 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24284__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18839__B2 _18792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25399_ _25411_/CLK _12711_/X HRESETn VGND VGND VPWR VPWR _12510_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15152_ _15143_/X _15146_/X _15152_/C _15152_/D VGND VGND VPWR VPWR _15162_/C sky130_fd_sc_hd__or4_4
X_12364_ _12364_/A VGND VGND VPWR VPWR _12364_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14103_ _14117_/C _14103_/B _25210_/Q VGND VGND VPWR VPWR _14103_/X sky130_fd_sc_hd__or3_4
XFILLER_5_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15083_ _15083_/A VGND VGND VPWR VPWR _15083_/Y sky130_fd_sc_hd__inv_2
X_19960_ _21929_/B _19957_/X _19622_/X _19957_/X VGND VGND VPWR VPWR _23545_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19498__A2_N _19495_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15522__B1 HADDR[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12295_ _12294_/Y _24838_/Q _12294_/Y _24838_/Q VGND VGND VPWR VPWR _12295_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22399__A1 _21493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14034_ _14032_/Y _14003_/B _14045_/A _14025_/D VGND VGND VPWR VPWR _14035_/A sky130_fd_sc_hd__or4_4
X_18911_ _23912_/Q VGND VGND VPWR VPWR _21755_/B sky130_fd_sc_hd__inv_2
XFILLER_10_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19891_ _19887_/Y _19890_/X _19612_/X _19890_/X VGND VGND VPWR VPWR _23572_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18842_ _16506_/A _24126_/Q _16506_/Y _18692_/A VGND VGND VPWR VPWR _18842_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25419__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15825__A1 _15824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15985_ _15788_/X _15857_/A _15768_/X _24738_/Q _15933_/A VGND VGND VPWR VPWR _15985_/X
+ sky130_fd_sc_hd__a32o_4
X_18773_ _18692_/B _18773_/B VGND VGND VPWR VPWR _18774_/A sky130_fd_sc_hd__or2_4
XANTENNA__13836__B1 _13835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25072__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14936_ _24997_/Q VGND VGND VPWR VPWR _15278_/A sky130_fd_sc_hd__inv_2
X_17724_ _17724_/A VGND VGND VPWR VPWR _17724_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25001__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14867_ _14811_/X _14866_/Y _24941_/Q _14811_/X VGND VGND VPWR VPWR _14867_/X sky130_fd_sc_hd__a2bb2o_4
X_17655_ _17657_/B VGND VGND VPWR VPWR _17656_/B sky130_fd_sc_hd__inv_2
XANTENNA__15589__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_37_0_HCLK clkbuf_6_18_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_75_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13818_ _21994_/A VGND VGND VPWR VPWR _18235_/A sky130_fd_sc_hd__buf_2
X_16606_ _24509_/Q VGND VGND VPWR VPWR _16606_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17586_ _24309_/Q _17586_/B VGND VGND VPWR VPWR _17588_/B sky130_fd_sc_hd__or2_4
X_14798_ _14869_/A _14798_/B _14870_/A _25031_/Q VGND VGND VPWR VPWR _14798_/X sky130_fd_sc_hd__or4_4
XFILLER_91_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16537_ _24535_/Q VGND VGND VPWR VPWR _16537_/Y sky130_fd_sc_hd__inv_2
X_19325_ _19311_/Y VGND VGND VPWR VPWR _19325_/X sky130_fd_sc_hd__buf_2
X_13749_ _13748_/C VGND VGND VPWR VPWR _13755_/A sky130_fd_sc_hd__inv_2
XANTENNA__20334__B1 _18267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12983__A _12983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16455__A _16725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16468_ _16465_/Y _16461_/X _16380_/X _16467_/X VGND VGND VPWR VPWR _16468_/X sky130_fd_sc_hd__a2bb2o_4
X_19256_ _19256_/A VGND VGND VPWR VPWR _19256_/X sky130_fd_sc_hd__buf_2
X_15419_ _15388_/B _15423_/A VGND VGND VPWR VPWR _15419_/Y sky130_fd_sc_hd__nand2_4
X_18207_ _18175_/A _23885_/Q VGND VGND VPWR VPWR _18208_/C sky130_fd_sc_hd__or2_4
X_19187_ _19187_/A VGND VGND VPWR VPWR _19187_/Y sky130_fd_sc_hd__inv_2
X_16399_ _15149_/Y _16394_/X _16398_/X _16394_/X VGND VGND VPWR VPWR _16399_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15761__B1 _15620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_6_0_HCLK clkbuf_3_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18138_ _18202_/A _18134_/X _18138_/C VGND VGND VPWR VPWR _18146_/B sky130_fd_sc_hd__or3_4
XFILLER_30_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18069_ _18217_/A _18065_/X _18069_/C VGND VGND VPWR VPWR _18078_/B sky130_fd_sc_hd__or3_4
X_20100_ _20098_/Y _20095_/X _20099_/X _20095_/X VGND VGND VPWR VPWR _20100_/X sky130_fd_sc_hd__a2bb2o_4
X_21080_ _21029_/X _21077_/X _21859_/C _21079_/X VGND VGND VPWR VPWR _21080_/X sky130_fd_sc_hd__a211o_4
XANTENNA__23936__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20031_ _23521_/Q VGND VGND VPWR VPWR _21920_/B sky130_fd_sc_hd__inv_2
XFILLER_112_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12223__A _25422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13827__B1 _11813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24770_ _23805_/CLK _15922_/X HRESETn VGND VGND VPWR VPWR _13540_/B sky130_fd_sc_hd__dfrtp_4
X_21982_ _21502_/X _21911_/X _21951_/X _21966_/Y _21981_/Y VGND VGND VPWR VPWR _21982_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_54_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23721_ _23887_/CLK _23721_/D VGND VGND VPWR VPWR _18073_/B sky130_fd_sc_hd__dfxtp_4
X_20933_ _20909_/X _20932_/X _24492_/Q _20913_/X VGND VGND VPWR VPWR _24055_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23652_ _23635_/CLK _23652_/D VGND VGND VPWR VPWR _19660_/A sky130_fd_sc_hd__dfxtp_4
X_20864_ _20913_/A VGND VGND VPWR VPWR _20864_/X sky130_fd_sc_hd__buf_2
XANTENNA__24795__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14989__A2_N _24448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22603_ _17744_/Y _22425_/A _12475_/A _22429_/A VGND VGND VPWR VPWR _22603_/X sky130_fd_sc_hd__o22a_4
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24724__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23583_ _24089_/CLK _19860_/X VGND VGND VPWR VPWR _19858_/A sky130_fd_sc_hd__dfxtp_4
X_20795_ _13136_/X VGND VGND VPWR VPWR _20800_/B sky130_fd_sc_hd__inv_2
XFILLER_74_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16365__A _24599_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21090__A1_N _21729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25322_ _25351_/CLK _25322_/D HRESETn VGND VGND VPWR VPWR _25322_/Q sky130_fd_sc_hd__dfrtp_4
X_22534_ _21303_/X VGND VGND VPWR VPWR _22534_/X sky130_fd_sc_hd__buf_2
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25253_ _25263_/CLK _25253_/D HRESETn VGND VGND VPWR VPWR _13544_/A sky130_fd_sc_hd__dfrtp_4
X_22465_ _22465_/A _23304_/B VGND VGND VPWR VPWR _22465_/X sky130_fd_sc_hd__or2_4
XFILLER_6_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22617__A2 _22614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12566__B1 _12565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24204_ _24288_/CLK _24204_/D HRESETn VGND VGND VPWR VPWR _17707_/A sky130_fd_sc_hd__dfrtp_4
X_21416_ _21416_/A VGND VGND VPWR VPWR _21416_/X sky130_fd_sc_hd__buf_2
X_25184_ _24942_/CLK _14234_/X HRESETn VGND VGND VPWR VPWR _25184_/Q sky130_fd_sc_hd__dfstp_4
X_22396_ _22394_/X _22395_/X _22396_/C VGND VGND VPWR VPWR _22396_/X sky130_fd_sc_hd__and3_4
X_24135_ _24136_/CLK _24135_/D HRESETn VGND VGND VPWR VPWR _18658_/A sky130_fd_sc_hd__dfrtp_4
X_21347_ _13468_/X _21345_/X _12054_/X _21346_/X VGND VGND VPWR VPWR _21347_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15709__A _15709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12080_ _12078_/Y _12074_/X _11842_/X _12079_/X VGND VGND VPWR VPWR _12080_/X sky130_fd_sc_hd__a2bb2o_4
X_24066_ _24069_/CLK _20524_/X HRESETn VGND VGND VPWR VPWR _24066_/Q sky130_fd_sc_hd__dfrtp_4
X_21278_ _21277_/Y VGND VGND VPWR VPWR _21278_/X sky130_fd_sc_hd__buf_2
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13229__A _13450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25512__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23017_ _23017_/A VGND VGND VPWR VPWR _23017_/Y sky130_fd_sc_hd__inv_2
X_20229_ _20228_/Y _20224_/X _19771_/X _20211_/Y VGND VGND VPWR VPWR _20229_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21446__A _17706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15770_ _12552_/Y _15763_/X _15477_/X _15763_/X VGND VGND VPWR VPWR _24844_/D sky130_fd_sc_hd__a2bb2o_4
X_12982_ _13042_/A VGND VGND VPWR VPWR _13038_/A sky130_fd_sc_hd__buf_2
XFILLER_92_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24968_ _24980_/CLK _15411_/X HRESETn VGND VGND VPWR VPWR _24968_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14491__B1 _14470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14721_ _14705_/A _14705_/B _21781_/A VGND VGND VPWR VPWR _14721_/X sky130_fd_sc_hd__and3_4
XFILLER_73_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11933_ _19618_/A VGND VGND VPWR VPWR _11933_/Y sky130_fd_sc_hd__inv_2
X_23919_ _24077_/CLK _23919_/D HRESETn VGND VGND VPWR VPWR _22306_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24899_ _24868_/CLK _24899_/D HRESETn VGND VGND VPWR VPWR _24899_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17440_ _17439_/X VGND VGND VPWR VPWR _21116_/A sky130_fd_sc_hd__buf_2
X_14652_ _17930_/A VGND VGND VPWR VPWR _17956_/A sky130_fd_sc_hd__buf_2
XFILLER_92_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11864_ _11864_/A VGND VGND VPWR VPWR _11864_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13603_ _25062_/Q VGND VGND VPWR VPWR _13610_/A sky130_fd_sc_hd__buf_2
X_17371_ _17371_/A VGND VGND VPWR VPWR _17372_/B sky130_fd_sc_hd__inv_2
XANTENNA__14794__A1 _13634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22708__C _21859_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14583_ _14581_/X _14557_/X _14582_/X _13770_/X _13568_/X VGND VGND VPWR VPWR _14583_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24465__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11795_ _11794_/X VGND VGND VPWR VPWR _11795_/X sky130_fd_sc_hd__buf_2
XANTENNA__19182__B1 _19136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16322_ _24615_/Q VGND VGND VPWR VPWR _16322_/Y sky130_fd_sc_hd__inv_2
X_19110_ _19109_/Y _19107_/X _18993_/X _19107_/X VGND VGND VPWR VPWR _19110_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13534_ _13534_/A VGND VGND VPWR VPWR _13534_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19041_ _19036_/Y _19040_/X _19018_/X _19040_/X VGND VGND VPWR VPWR _19041_/X sky130_fd_sc_hd__a2bb2o_4
X_16253_ _22154_/A VGND VGND VPWR VPWR _16253_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13465_ _23343_/A VGND VGND VPWR VPWR _13465_/Y sky130_fd_sc_hd__inv_2
X_15204_ _15198_/A _15204_/B _15203_/X VGND VGND VPWR VPWR _15204_/X sky130_fd_sc_hd__and3_4
X_12416_ _12277_/B _12415_/X VGND VGND VPWR VPWR _12419_/B sky130_fd_sc_hd__or2_4
XFILLER_103_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16184_ _16184_/A VGND VGND VPWR VPWR _16459_/B sky130_fd_sc_hd__buf_2
XFILLER_51_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13396_ _13428_/A _13396_/B _13395_/X VGND VGND VPWR VPWR _13396_/X sky130_fd_sc_hd__and3_4
XFILLER_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17818__B _17758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15135_ _24986_/Q VGND VGND VPWR VPWR _15135_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12347_ _25334_/Q VGND VGND VPWR VPWR _12347_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12762__A2_N _24772_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15066_ _14960_/Y _14949_/Y _15065_/Y _15212_/A VGND VGND VPWR VPWR _15068_/C sky130_fd_sc_hd__or4_4
X_19943_ _19943_/A VGND VGND VPWR VPWR _19943_/X sky130_fd_sc_hd__buf_2
X_12278_ _12475_/A _12278_/B _12278_/C _12196_/Y VGND VGND VPWR VPWR _12278_/X sky130_fd_sc_hd__or4_4
XANTENNA__13784__D _13784_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22740__A _24750_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14017_ _14002_/X VGND VGND VPWR VPWR _14017_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25253__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19874_ _19872_/Y _19868_/X _19618_/X _19873_/X VGND VGND VPWR VPWR _23578_/D sky130_fd_sc_hd__a2bb2o_4
X_18825_ _16501_/Y _18767_/A _16501_/Y _18767_/A VGND VGND VPWR VPWR _18825_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12978__A _25355_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18756_ _18753_/C _18756_/B VGND VGND VPWR VPWR _18757_/B sky130_fd_sc_hd__or2_4
X_15968_ _15966_/X _15935_/X HWDATA[16] _24751_/Q _15967_/X VGND VGND VPWR VPWR _15968_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14482__B1 _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17707_ _17707_/A VGND VGND VPWR VPWR _17708_/A sky130_fd_sc_hd__buf_2
X_14919_ _14919_/A VGND VGND VPWR VPWR _14919_/Y sky130_fd_sc_hd__inv_2
X_15899_ _12785_/Y _15896_/X _15756_/X _15896_/X VGND VGND VPWR VPWR _15899_/X sky130_fd_sc_hd__a2bb2o_4
X_18687_ _24128_/Q VGND VGND VPWR VPWR _18768_/A sky130_fd_sc_hd__inv_2
XFILLER_110_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17638_ _17567_/A _17642_/B _17637_/Y VGND VGND VPWR VPWR _17638_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14234__B1 _13800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22187__A _22153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17569_ _17630_/A _17541_/Y _17568_/X VGND VGND VPWR VPWR _17569_/X sky130_fd_sc_hd__or3_4
XANTENNA__22847__A2 _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16185__A _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19308_ _19306_/Y _19302_/X _19307_/X _19287_/Y VGND VGND VPWR VPWR _19308_/X sky130_fd_sc_hd__a2bb2o_4
X_20580_ _14421_/Y _20556_/A _20546_/X _20579_/X VGND VGND VPWR VPWR _20580_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24135__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_124_0_HCLK clkbuf_7_62_0_HCLK/X VGND VGND VPWR VPWR _24465_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22915__A _22915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20322__A3 _13835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_187_0_HCLK clkbuf_7_93_0_HCLK/X VGND VGND VPWR VPWR _23550_/CLK sky130_fd_sc_hd__clkbuf_1
X_19239_ _13436_/B VGND VGND VPWR VPWR _19239_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15734__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22250_ _22246_/A _22250_/B VGND VGND VPWR VPWR _22250_/X sky130_fd_sc_hd__or2_4
X_21201_ _13791_/X _21198_/X _21200_/X _23342_/A _21996_/A VGND VGND VPWR VPWR _21201_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_69_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22181_ _22181_/A _21220_/A VGND VGND VPWR VPWR _22186_/B sky130_fd_sc_hd__or2_4
XANTENNA__15529__A _15535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14433__A _14433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21132_ _21014_/A _21131_/X VGND VGND VPWR VPWR _21132_/Y sky130_fd_sc_hd__nor2_4
X_21063_ _21062_/Y VGND VGND VPWR VPWR _21064_/A sky130_fd_sc_hd__buf_2
XFILLER_8_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20014_ _20014_/A VGND VGND VPWR VPWR _20014_/X sky130_fd_sc_hd__buf_2
XFILLER_115_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12888__A _12841_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24822_ _24018_/CLK _15820_/X HRESETn VGND VGND VPWR VPWR _24822_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24976__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24753_ _24759_/CLK _15963_/X HRESETn VGND VGND VPWR VPWR _22853_/A sky130_fd_sc_hd__dfrtp_4
X_21965_ _21816_/B _21952_/X _21956_/Y _13784_/D _21964_/X VGND VGND VPWR VPWR _21965_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24905__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _23711_/CLK _23704_/D VGND VGND VPWR VPWR _23704_/Q sky130_fd_sc_hd__dfxtp_4
X_20916_ _24051_/Q _20911_/X _20915_/Y VGND VGND VPWR VPWR _20916_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14225__B1 _13835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21713__B _21713_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24684_ _24689_/CLK _16127_/X HRESETn VGND VGND VPWR VPWR _22774_/A sky130_fd_sc_hd__dfrtp_4
X_21896_ _14689_/A _20156_/Y VGND VGND VPWR VPWR _21896_/X sky130_fd_sc_hd__or2_4
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_20_0_HCLK clkbuf_7_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_20_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22299__B1 _22885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _23635_/CLK _23635_/D VGND VGND VPWR VPWR _13247_/B sky130_fd_sc_hd__dfxtp_4
X_20847_ _13659_/A _13659_/B VGND VGND VPWR VPWR _20847_/X sky130_fd_sc_hd__or2_4
XANTENNA__15973__B1 _24747_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_83_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_83_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23566_ _23550_/CLK _19905_/X VGND VGND VPWR VPWR _23566_/Q sky130_fd_sc_hd__dfxtp_4
X_20778_ _20770_/X _20777_/Y _15583_/A _20774_/X VGND VGND VPWR VPWR _20778_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25305_ _25305_/CLK _25305_/D HRESETn VGND VGND VPWR VPWR _25305_/Q sky130_fd_sc_hd__dfrtp_4
X_22517_ _22514_/X _22782_/A VGND VGND VPWR VPWR _22518_/D sky130_fd_sc_hd__nor2_4
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23497_ _23496_/CLK _20090_/X VGND VGND VPWR VPWR _23497_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ _13453_/A _13250_/B _13249_/X VGND VGND VPWR VPWR _13255_/B sky130_fd_sc_hd__and3_4
X_25236_ _25172_/CLK _25236_/D HRESETn VGND VGND VPWR VPWR _22111_/A sky130_fd_sc_hd__dfrtp_4
X_22448_ _16249_/Y _22444_/X _15099_/Y _22441_/X VGND VGND VPWR VPWR _22449_/B sky130_fd_sc_hd__o22a_4
XFILLER_100_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23263__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20345__A _20339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12201_ _12199_/A _22853_/A _12199_/Y _12200_/Y VGND VGND VPWR VPWR _12201_/X sky130_fd_sc_hd__o22a_4
X_13181_ _13168_/A _13179_/X _13180_/X VGND VGND VPWR VPWR _13181_/X sky130_fd_sc_hd__and3_4
X_25167_ _25461_/CLK _25167_/D HRESETn VGND VGND VPWR VPWR _25167_/Q sky130_fd_sc_hd__dfrtp_4
X_22379_ _21767_/X _22378_/X _14714_/X VGND VGND VPWR VPWR _22379_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_89_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12132_ _12126_/B VGND VGND VPWR VPWR _12132_/Y sky130_fd_sc_hd__inv_2
X_24118_ _24117_/CLK _24118_/D HRESETn VGND VGND VPWR VPWR _18809_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16150__B1 _16057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23015__A2 _22824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25098_ _25098_/CLK _25098_/D HRESETn VGND VGND VPWR VPWR _20441_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22223__B1 _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12063_ _12063_/A VGND VGND VPWR VPWR _12063_/Y sky130_fd_sc_hd__inv_2
X_16940_ _16156_/Y _17745_/A _23219_/A _16939_/Y VGND VGND VPWR VPWR _16940_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24049_ _24049_/CLK _20908_/X HRESETn VGND VGND VPWR VPWR _24049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16871_ _19787_/A VGND VGND VPWR VPWR _16871_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18610_ _18610_/A VGND VGND VPWR VPWR _18610_/Y sky130_fd_sc_hd__inv_2
X_15822_ _15816_/X _15819_/X _11809_/A _24820_/Q _15817_/X VGND VGND VPWR VPWR _15822_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17650__B1 _17601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19590_ _22220_/A VGND VGND VPWR VPWR _19590_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15753_ _15749_/X _15742_/X _15752_/X _24853_/Q _15711_/A VGND VGND VPWR VPWR _15753_/X
+ sky130_fd_sc_hd__a32o_4
X_18541_ _18541_/A _18541_/B _18540_/Y VGND VGND VPWR VPWR _24162_/D sky130_fd_sc_hd__and3_4
X_12965_ _12959_/B VGND VGND VPWR VPWR _12966_/B sky130_fd_sc_hd__inv_2
XANTENNA__24646__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22719__B _22693_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11916_ _11916_/A _11916_/B VGND VGND VPWR VPWR _11916_/X sky130_fd_sc_hd__and2_4
X_14704_ _14675_/X VGND VGND VPWR VPWR _14705_/B sky130_fd_sc_hd__inv_2
X_15684_ _15684_/A VGND VGND VPWR VPWR _15685_/A sky130_fd_sc_hd__inv_2
X_18472_ _18472_/A _18418_/Y _18471_/Y _18566_/A VGND VGND VPWR VPWR _18476_/B sky130_fd_sc_hd__or4_4
X_12896_ _12896_/A _12896_/B VGND VGND VPWR VPWR _12897_/C sky130_fd_sc_hd__or2_4
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14635_ _14634_/Y _14622_/Y _14632_/A _14622_/A VGND VGND VPWR VPWR _14635_/X sky130_fd_sc_hd__o22a_4
X_17423_ _17423_/A VGND VGND VPWR VPWR _17423_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11847_ _16355_/A VGND VGND VPWR VPWR _11847_/X sky130_fd_sc_hd__buf_2
XFILLER_18_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13422__A _13454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14566_ _14559_/Y _14596_/B VGND VGND VPWR VPWR _14567_/B sky130_fd_sc_hd__or2_4
X_17354_ _17370_/A _17354_/B _17354_/C VGND VGND VPWR VPWR _24339_/D sky130_fd_sc_hd__and3_4
XFILLER_57_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11778_ HWDATA[21] VGND VGND VPWR VPWR _11778_/X sky130_fd_sc_hd__buf_2
XFILLER_105_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13517_ _25294_/Q VGND VGND VPWR VPWR _13517_/Y sky130_fd_sc_hd__inv_2
X_16305_ _23039_/A VGND VGND VPWR VPWR _16305_/Y sky130_fd_sc_hd__inv_2
X_17285_ _17178_/Y _17283_/A VGND VGND VPWR VPWR _17285_/X sky130_fd_sc_hd__or2_4
X_14497_ _14541_/A _14495_/X _14496_/X VGND VGND VPWR VPWR _14497_/X sky130_fd_sc_hd__o21a_4
XFILLER_118_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16733__A _16733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18662__A1_N _16547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16236_ _16234_/Y _16232_/X _16235_/X _16232_/X VGND VGND VPWR VPWR _24647_/D sky130_fd_sc_hd__a2bb2o_4
X_19024_ _19022_/Y _19016_/X _18997_/X _19023_/X VGND VGND VPWR VPWR _23874_/D sky130_fd_sc_hd__a2bb2o_4
X_13448_ _13310_/A _23645_/Q VGND VGND VPWR VPWR _13448_/X sky130_fd_sc_hd__or2_4
X_16167_ _14781_/A _14764_/Y VGND VGND VPWR VPWR _16167_/X sky130_fd_sc_hd__and2_4
XANTENNA__25434__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13379_ _13379_/A _13379_/B VGND VGND VPWR VPWR _13379_/X sky130_fd_sc_hd__or2_4
XANTENNA__13795__C _13784_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15118_ _24585_/Q VGND VGND VPWR VPWR _15118_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16098_ _23187_/A VGND VGND VPWR VPWR _16098_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16141__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23006__A2 _22393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15049_ _14888_/Y _24464_/Q _14888_/Y _24464_/Q VGND VGND VPWR VPWR _15049_/X sky130_fd_sc_hd__a2bb2o_4
X_19926_ _19925_/Y _19923_/X _19797_/X _19923_/X VGND VGND VPWR VPWR _19926_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17564__A _24294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23285__B _23226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21086__A _24599_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19857_ _21764_/B _19852_/X _19790_/X _19852_/X VGND VGND VPWR VPWR _19857_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18600__A1_N _16541_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18808_ _18786_/D VGND VGND VPWR VPWR _18809_/B sky130_fd_sc_hd__inv_2
XFILLER_56_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19788_ _21881_/B _19784_/X _19787_/X _19784_/X VGND VGND VPWR VPWR _19788_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21814__A _21681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18739_ _18693_/X _18703_/X _18658_/Y VGND VGND VPWR VPWR _18740_/C sky130_fd_sc_hd__o21a_4
XFILLER_97_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24387__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21750_ _21609_/A _21750_/B _21749_/X VGND VGND VPWR VPWR _21750_/X sky130_fd_sc_hd__and3_4
XFILLER_3_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24316__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18615__A1_N _16622_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24547__D _16507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20701_ _15625_/Y _20698_/X _20686_/X _20700_/X VGND VGND VPWR VPWR _20702_/A sky130_fd_sc_hd__o22a_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21681_ _21681_/A _21672_/X _21681_/C VGND VGND VPWR VPWR _21681_/X sky130_fd_sc_hd__or3_4
XANTENNA__14428__A _25126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23420_ _23396_/CLK _23420_/D VGND VGND VPWR VPWR _23420_/Q sky130_fd_sc_hd__dfxtp_4
X_20632_ _20632_/A VGND VGND VPWR VPWR _20632_/Y sky130_fd_sc_hd__inv_2
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15970__A3 _11800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23351_ VGND VGND VPWR VPWR _23351_/HI scl_o_S5 sky130_fd_sc_hd__conb_1
X_20563_ _20566_/B _20561_/Y _20571_/C VGND VGND VPWR VPWR _20563_/X sky130_fd_sc_hd__and3_4
XFILLER_123_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22302_ _22302_/A _22316_/B VGND VGND VPWR VPWR _22302_/Y sky130_fd_sc_hd__nor2_4
X_23282_ _12266_/Y _21524_/X _24275_/Q _22483_/X VGND VGND VPWR VPWR _23282_/X sky130_fd_sc_hd__a2bb2o_4
X_20494_ _20494_/A _20493_/X VGND VGND VPWR VPWR _20494_/X sky130_fd_sc_hd__or2_4
XANTENNA__23951__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25021_ _25024_/CLK _15191_/Y HRESETn VGND VGND VPWR VPWR _25021_/Q sky130_fd_sc_hd__dfrtp_4
X_22233_ _17720_/X _22228_/X _22232_/X VGND VGND VPWR VPWR _22233_/X sky130_fd_sc_hd__or3_4
XANTENNA__22453__B1 _13813_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11787__A _25525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11744__B2 _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25104__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22164_ _14478_/Y _14257_/A _25095_/Q _22172_/B VGND VGND VPWR VPWR _22164_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16132__B1 _11804_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21115_ _21101_/Y _21103_/X _21106_/X _21114_/X VGND VGND VPWR VPWR _21272_/A sky130_fd_sc_hd__a211o_4
XFILLER_132_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17474__A _17474_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22095_ _14441_/Y _21352_/A _14458_/Y _17415_/A VGND VGND VPWR VPWR _22095_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22756__B2 _22755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20789__A1_N _20770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21046_ _21015_/A VGND VGND VPWR VPWR _21306_/A sky130_fd_sc_hd__buf_2
XFILLER_87_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17632__B1 _17601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24805_ _24025_/CLK _24805_/D HRESETn VGND VGND VPWR VPWR _12604_/A sky130_fd_sc_hd__dfrtp_4
X_22997_ _22997_/A VGND VGND VPWR VPWR _22997_/X sky130_fd_sc_hd__buf_2
XANTENNA__19385__B1 _19294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22539__B _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12750_ _12749_/Y _24797_/Q _12749_/Y _24797_/Q VGND VGND VPWR VPWR _12750_/X sky130_fd_sc_hd__a2bb2o_4
X_24736_ _25374_/CLK _24736_/D HRESETn VGND VGND VPWR VPWR _21433_/A sky130_fd_sc_hd__dfrtp_4
X_21948_ _21681_/A _21940_/X _21948_/C VGND VGND VPWR VPWR _21948_/X sky130_fd_sc_hd__or3_4
XANTENNA__24057__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11701_/A _11701_/B _11700_/X VGND VGND VPWR VPWR _17445_/C sky130_fd_sc_hd__or3_4
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12681_/A _12684_/B VGND VGND VPWR VPWR _12682_/C sky130_fd_sc_hd__nand2_4
XANTENNA__15946__B1 _15944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24667_ _23467_/CLK _16177_/X HRESETn VGND VGND VPWR VPWR _13738_/A sky130_fd_sc_hd__dfrtp_4
X_21879_ _14693_/A _21879_/B _21878_/X VGND VGND VPWR VPWR _21879_/X sky130_fd_sc_hd__and3_4
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14416_/Y _14409_/X _14418_/X _14419_/X VGND VGND VPWR VPWR _25130_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _23618_/CLK _23618_/D VGND VGND VPWR VPWR _19757_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24598_ _24984_/CLK _24598_/D HRESETn VGND VGND VPWR VPWR _24598_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14351_ _14348_/Y VGND VGND VPWR VPWR _14351_/X sky130_fd_sc_hd__buf_2
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22692__B1 _22783_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23549_ _24309_/CLK _19948_/X VGND VGND VPWR VPWR _23549_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16553__A _24530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _13225_/A VGND VGND VPWR VPWR _13303_/A sky130_fd_sc_hd__buf_2
X_17070_ _17060_/B VGND VGND VPWR VPWR _17071_/B sky130_fd_sc_hd__inv_2
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _20488_/A VGND VGND VPWR VPWR _14282_/X sky130_fd_sc_hd__buf_2
XFILLER_52_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_170_0_HCLK clkbuf_7_85_0_HCLK/X VGND VGND VPWR VPWR _24923_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16021_ _24724_/Q VGND VGND VPWR VPWR _16021_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13233_ _13233_/A VGND VGND VPWR VPWR _13386_/A sky130_fd_sc_hd__buf_2
XANTENNA__15169__A _14888_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_27_0_HCLK clkbuf_8_27_0_HCLK/A VGND VGND VPWR VPWR _25284_/CLK sky130_fd_sc_hd__clkbuf_1
X_25219_ _25219_/CLK _14085_/X HRESETn VGND VGND VPWR VPWR _25219_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13164_ _13186_/A _23636_/Q VGND VGND VPWR VPWR _13164_/X sky130_fd_sc_hd__or2_4
XANTENNA__16123__B1 _15964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12115_ _12113_/Y _12114_/X _11847_/X _12114_/X VGND VGND VPWR VPWR _12115_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17384__A _17242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13095_ _13076_/A _13092_/B _13095_/C VGND VGND VPWR VPWR _13095_/X sky130_fd_sc_hd__and3_4
X_17972_ _13610_/A VGND VGND VPWR VPWR _17996_/A sky130_fd_sc_hd__buf_2
XFILLER_78_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24898__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19711_ _23634_/Q VGND VGND VPWR VPWR _19711_/Y sky130_fd_sc_hd__inv_2
X_12046_ _23344_/A VGND VGND VPWR VPWR _12046_/Y sky130_fd_sc_hd__inv_2
X_16923_ _16895_/X _16904_/X _16913_/X _16922_/X VGND VGND VPWR VPWR _16953_/A sky130_fd_sc_hd__or4_4
XANTENNA__18415__A2 _18414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24827__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19642_ _19642_/A VGND VGND VPWR VPWR _19642_/X sky130_fd_sc_hd__buf_2
XANTENNA__13417__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16854_ _14944_/Y _16796_/X _16717_/X _16796_/X VGND VGND VPWR VPWR _24402_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15805_ _15781_/X _15795_/X _15725_/X _24832_/Q _15793_/X VGND VGND VPWR VPWR _15805_/X
+ sky130_fd_sc_hd__a32o_4
X_19573_ _23679_/Q VGND VGND VPWR VPWR _19573_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24480__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13997_ _13997_/A VGND VGND VPWR VPWR _13997_/X sky130_fd_sc_hd__buf_2
X_16785_ _16785_/A VGND VGND VPWR VPWR _16785_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16728__A _16728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18524_ _18524_/A _18523_/X VGND VGND VPWR VPWR _18525_/A sky130_fd_sc_hd__or2_4
XFILLER_0_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15632__A _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12948_ _12964_/A _12946_/X _12947_/X VGND VGND VPWR VPWR _25366_/D sky130_fd_sc_hd__and3_4
X_15736_ _12533_/Y _15732_/X _11784_/X _15735_/X VGND VGND VPWR VPWR _24861_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18455_ _18455_/A VGND VGND VPWR VPWR _18482_/A sky130_fd_sc_hd__inv_2
XANTENNA__15351__B _15336_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12879_ _12747_/A _12879_/B VGND VGND VPWR VPWR _12879_/X sky130_fd_sc_hd__or2_4
X_15667_ _15667_/A VGND VGND VPWR VPWR _15668_/A sky130_fd_sc_hd__buf_2
XFILLER_33_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13152__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17406_ _17387_/X _17401_/X _20992_/B _24326_/Q _17404_/X VGND VGND VPWR VPWR _17406_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14618_ _14615_/Y _13638_/X _14617_/Y VGND VGND VPWR VPWR _14630_/B sky130_fd_sc_hd__o21ai_4
X_15598_ _22787_/A _15593_/X _11796_/X _15593_/X VGND VGND VPWR VPWR _15598_/X sky130_fd_sc_hd__a2bb2o_4
X_18386_ _24179_/Q VGND VGND VPWR VPWR _18386_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12215__A2 _22892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14549_ _14542_/X _14548_/Y sda_oen_o_S4 _14542_/X VGND VGND VPWR VPWR _25087_/D
+ sky130_fd_sc_hd__a2bb2o_4
X_17337_ _17249_/Y _17336_/X VGND VGND VPWR VPWR _17337_/X sky130_fd_sc_hd__or2_4
XFILLER_18_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16463__A _24564_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17268_ _17260_/B _17267_/X VGND VGND VPWR VPWR _17269_/C sky130_fd_sc_hd__or2_4
XFILLER_105_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16362__B1 _15986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19007_ _19007_/A VGND VGND VPWR VPWR _19007_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16219_ _22878_/A VGND VGND VPWR VPWR _16219_/Y sky130_fd_sc_hd__inv_2
X_17199_ _17199_/A VGND VGND VPWR VPWR _17199_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19300__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16114__B1 _15955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19909_ _13755_/A _13752_/X _20043_/A _13762_/A VGND VGND VPWR VPWR _19909_/X sky130_fd_sc_hd__or4_4
XANTENNA__24568__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13327__A _13233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17614__B1 _17590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22920_ _23056_/A _22919_/Y VGND VGND VPWR VPWR _22920_/Y sky130_fd_sc_hd__nor2_4
XFILLER_25_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12231__A _21433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22851_ _22842_/Y _22849_/Y _22850_/X VGND VGND VPWR VPWR _22851_/X sky130_fd_sc_hd__o21a_4
XFILLER_44_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14979__B2 _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19367__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21802_ _21649_/A _21800_/X _21801_/X VGND VGND VPWR VPWR _21802_/X sky130_fd_sc_hd__and3_4
XANTENNA__24150__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22782_ _22782_/A VGND VGND VPWR VPWR _23054_/A sky130_fd_sc_hd__buf_2
XFILLER_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12593__A2_N _24872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24521_ _24555_/CLK _24521_/D HRESETn VGND VGND VPWR VPWR _24521_/Q sky130_fd_sc_hd__dfrtp_4
X_21733_ _16850_/Y _15708_/A _21316_/A _21732_/X VGND VGND VPWR VPWR _21733_/X sky130_fd_sc_hd__o22a_4
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24452_ _25024_/CLK _16754_/X HRESETn VGND VGND VPWR VPWR _24452_/Q sky130_fd_sc_hd__dfrtp_4
X_21664_ _21664_/A _20372_/Y VGND VGND VPWR VPWR _21664_/X sky130_fd_sc_hd__or2_4
XANTENNA__22269__A3 _21290_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25132__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23403_ _23580_/CLK _20341_/X VGND VGND VPWR VPWR _20337_/A sky130_fd_sc_hd__dfxtp_4
X_20615_ _20620_/B _20615_/B _20611_/C VGND VGND VPWR VPWR _20615_/X sky130_fd_sc_hd__and3_4
XFILLER_138_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25356__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22674__B1 _22613_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24383_ _24383_/CLK _24383_/D HRESETn VGND VGND VPWR VPWR _17085_/A sky130_fd_sc_hd__dfrtp_4
X_21595_ _21595_/A VGND VGND VPWR VPWR _21596_/A sky130_fd_sc_hd__buf_2
XFILLER_137_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16373__A _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23334_ _13802_/Y _25057_/Q _21366_/A _13598_/C VGND VGND VPWR VPWR _23334_/X sky130_fd_sc_hd__o22a_4
X_20546_ _14381_/A VGND VGND VPWR VPWR _20546_/X sky130_fd_sc_hd__buf_2
XANTENNA__16353__B1 _16064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_243_0_HCLK clkbuf_8_243_0_HCLK/A VGND VGND VPWR VPWR _24865_/CLK sky130_fd_sc_hd__clkbuf_1
X_23265_ _21438_/X _23263_/X _22684_/X _23264_/X VGND VGND VPWR VPWR _23265_/X sky130_fd_sc_hd__o22a_4
X_20477_ _20506_/A _20473_/X _20486_/B VGND VGND VPWR VPWR _20502_/A sky130_fd_sc_hd__o21a_4
X_25004_ _25001_/CLK _15263_/X HRESETn VGND VGND VPWR VPWR _25004_/Q sky130_fd_sc_hd__dfrtp_4
X_22216_ _21622_/A _22216_/B VGND VGND VPWR VPWR _22216_/X sky130_fd_sc_hd__or2_4
XFILLER_134_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23196_ _23119_/X _23194_/X _23121_/X _23195_/X VGND VGND VPWR VPWR _23197_/B sky130_fd_sc_hd__o22a_4
XFILLER_117_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22147_ _21098_/X _22140_/X _22143_/X _22146_/X VGND VGND VPWR VPWR _22148_/B sky130_fd_sc_hd__a211o_4
XFILLER_117_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14206__A1_N _14205_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24991__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22078_ _21377_/A VGND VGND VPWR VPWR _22078_/X sky130_fd_sc_hd__buf_2
XFILLER_0_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24920__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13920_ _13920_/A VGND VGND VPWR VPWR _13920_/X sky130_fd_sc_hd__buf_2
X_21029_ _21112_/B VGND VGND VPWR VPWR _21029_/X sky130_fd_sc_hd__buf_2
XFILLER_120_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24238__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_12_0_HCLK_A clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13851_ _13851_/A _20466_/B _13850_/Y VGND VGND VPWR VPWR _13851_/X sky130_fd_sc_hd__or3_4
XANTENNA__21454__A _21454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12802_ _12849_/B VGND VGND VPWR VPWR _12924_/A sky130_fd_sc_hd__buf_2
X_13782_ _13782_/A VGND VGND VPWR VPWR _13782_/X sky130_fd_sc_hd__buf_2
X_16570_ _16558_/A VGND VGND VPWR VPWR _16570_/X sky130_fd_sc_hd__buf_2
XFILLER_16_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12733_ _12729_/A _12737_/A VGND VGND VPWR VPWR _12734_/B sky130_fd_sc_hd__nand2_4
X_15521_ _11730_/B VGND VGND VPWR VPWR _15521_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15171__B _15171_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24719_ _24345_/CLK _16036_/X HRESETn VGND VGND VPWR VPWR _16033_/A sky130_fd_sc_hd__dfrtp_4
X_15452_ _15452_/A VGND VGND VPWR VPWR _15452_/X sky130_fd_sc_hd__buf_2
X_18240_ _11697_/Y _18233_/X _15747_/X _18233_/X VGND VGND VPWR VPWR _24226_/D sky130_fd_sc_hd__a2bb2o_4
X_12664_ _12664_/A VGND VGND VPWR VPWR _12686_/A sky130_fd_sc_hd__buf_2
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15934__A3 _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _16359_/A VGND VGND VPWR VPWR _14403_/X sky130_fd_sc_hd__buf_2
XFILLER_54_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25097__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_53_0_HCLK clkbuf_6_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15383_ _15133_/Y _15380_/X VGND VGND VPWR VPWR _15384_/C sky130_fd_sc_hd__or2_4
X_18171_ _18024_/A _18171_/B VGND VGND VPWR VPWR _18171_/X sky130_fd_sc_hd__or2_4
XANTENNA__22665__B1 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _12595_/A VGND VGND VPWR VPWR _12595_/Y sky130_fd_sc_hd__inv_2
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14334_ _18370_/B _14333_/X _14325_/X VGND VGND VPWR VPWR _25154_/D sky130_fd_sc_hd__a21o_4
X_17122_ _17036_/A _17121_/Y VGND VGND VPWR VPWR _17122_/X sky130_fd_sc_hd__or2_4
XFILLER_89_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11956__B2 _11947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25026__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16344__B1 _16143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17053_ _24391_/Q _17053_/B VGND VGND VPWR VPWR _17054_/C sky130_fd_sc_hd__nand2_4
XFILLER_13_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14265_ _14263_/Y _14259_/X _13840_/X _14264_/X VGND VGND VPWR VPWR _25177_/D sky130_fd_sc_hd__a2bb2o_4
X_16004_ _16001_/Y _15997_/X _15940_/X _16003_/X VGND VGND VPWR VPWR _16004_/X sky130_fd_sc_hd__a2bb2o_4
X_13216_ _13454_/A _13207_/X _13215_/X VGND VGND VPWR VPWR _13216_/X sky130_fd_sc_hd__or3_4
XFILLER_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14196_ _20467_/A _20476_/A VGND VGND VPWR VPWR _14196_/X sky130_fd_sc_hd__or2_4
XFILLER_83_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23090__B1 _11766_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13147_ _13234_/A VGND VGND VPWR VPWR _13251_/A sky130_fd_sc_hd__buf_2
XANTENNA__15627__A _16528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21640__A1 _21636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21640__B2 _18261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18003__A _18010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13078_ _13077_/X VGND VGND VPWR VPWR _25334_/D sky130_fd_sc_hd__inv_2
X_17955_ _17955_/A _23724_/Q VGND VGND VPWR VPWR _17957_/B sky130_fd_sc_hd__or2_4
XFILLER_61_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24661__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12029_ _12034_/A VGND VGND VPWR VPWR _12029_/X sky130_fd_sc_hd__buf_2
X_16906_ _22865_/A _24263_/Q _16120_/Y _17758_/A VGND VGND VPWR VPWR _16906_/X sky130_fd_sc_hd__o22a_4
X_17886_ _17737_/X _17848_/B _17885_/X VGND VGND VPWR VPWR _24245_/D sky130_fd_sc_hd__and3_4
XFILLER_93_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19625_ _11948_/A VGND VGND VPWR VPWR _19625_/X sky130_fd_sc_hd__buf_2
X_16837_ _16840_/A VGND VGND VPWR VPWR _16837_/X sky130_fd_sc_hd__buf_2
XFILLER_38_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12986__A _12299_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19556_ _19555_/Y _19552_/X _19462_/X _19552_/X VGND VGND VPWR VPWR _23686_/D sky130_fd_sc_hd__a2bb2o_4
X_16768_ _16767_/Y _16764_/X _15750_/X _16764_/X VGND VGND VPWR VPWR _16768_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21156__B1 _21314_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18507_ _18507_/A VGND VGND VPWR VPWR _24171_/D sky130_fd_sc_hd__inv_2
X_15719_ _12546_/Y _15718_/X _11749_/X _15718_/X VGND VGND VPWR VPWR _15719_/X sky130_fd_sc_hd__a2bb2o_4
X_19487_ _23709_/Q VGND VGND VPWR VPWR _19487_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20903__B1 _20845_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16699_ _16699_/A VGND VGND VPWR VPWR _16699_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18438_ _18438_/A VGND VGND VPWR VPWR _18456_/A sky130_fd_sc_hd__inv_2
XANTENNA__17289__A _17289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18369_ _18369_/A VGND VGND VPWR VPWR _18369_/Y sky130_fd_sc_hd__inv_2
X_20400_ _20399_/Y VGND VGND VPWR VPWR _20400_/X sky130_fd_sc_hd__buf_2
XANTENNA__13610__A _13610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21380_ _14679_/A VGND VGND VPWR VPWR _21381_/A sky130_fd_sc_hd__buf_2
XANTENNA__16335__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22923__A _22923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20331_ _20331_/A VGND VGND VPWR VPWR _20331_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22408__B1 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_10_0_HCLK clkbuf_7_5_0_HCLK/X VGND VGND VPWR VPWR _23516_/CLK sky130_fd_sc_hd__clkbuf_1
X_23050_ _23048_/X _23049_/X _23117_/C VGND VGND VPWR VPWR _23050_/X sky130_fd_sc_hd__or3_4
X_20262_ _21903_/B _20259_/X _19787_/A _20259_/X VGND VGND VPWR VPWR _23433_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22423__A3 _22422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24749__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22001_ _21194_/A VGND VGND VPWR VPWR _22247_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_73_0_HCLK clkbuf_8_73_0_HCLK/A VGND VGND VPWR VPWR _24945_/CLK sky130_fd_sc_hd__clkbuf_1
X_20193_ _23459_/Q VGND VGND VPWR VPWR _22216_/B sky130_fd_sc_hd__inv_2
XFILLER_89_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14441__A _25122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23952_ _24077_/CLK _23952_/D HRESETn VGND VGND VPWR VPWR _23952_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24331__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22903_ _15791_/A _22902_/X _22485_/X _25526_/Q _22775_/X VGND VGND VPWR VPWR _22903_/X
+ sky130_fd_sc_hd__a32o_4
X_23883_ _23884_/CLK _18994_/X VGND VGND VPWR VPWR _18991_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_57_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15074__B1 _15073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12896__A _12896_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22089__B _23082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22834_ _22923_/A VGND VGND VPWR VPWR _22834_/X sky130_fd_sc_hd__buf_2
XFILLER_25_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21698__A1 _16640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21698__B2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25537__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22765_ _24788_/Q _22472_/B VGND VGND VPWR VPWR _22765_/X sky130_fd_sc_hd__or2_4
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19760__B1 _19758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24504_ _24541_/CLK _24504_/D HRESETn VGND VGND VPWR VPWR _16618_/A sky130_fd_sc_hd__dfrtp_4
X_21716_ _21716_/A VGND VGND VPWR VPWR _21716_/Y sky130_fd_sc_hd__inv_2
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25484_ _23689_/CLK _11986_/X HRESETn VGND VGND VPWR VPWR _11654_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22696_ _24415_/Q _22406_/B _15667_/A _22695_/X VGND VGND VPWR VPWR _22696_/X sky130_fd_sc_hd__a211o_4
XANTENNA__20618__A _14807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24435_ _24435_/CLK _16789_/X HRESETn VGND VGND VPWR VPWR _24435_/Q sky130_fd_sc_hd__dfrtp_4
X_21647_ _21449_/A _19506_/Y VGND VGND VPWR VPWR _21647_/X sky130_fd_sc_hd__or2_4
XFILLER_36_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12380_ _12373_/X _12380_/B _12380_/C _12379_/X VGND VGND VPWR VPWR _12380_/X sky130_fd_sc_hd__or4_4
XANTENNA__16326__B1 _16325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24366_ _24362_/CLK _17148_/X HRESETn VGND VGND VPWR VPWR _16960_/A sky130_fd_sc_hd__dfrtp_4
X_21578_ _15668_/X _21578_/B VGND VGND VPWR VPWR _21578_/Y sky130_fd_sc_hd__nor2_4
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23317_ _23317_/A _16795_/A VGND VGND VPWR VPWR _23317_/Y sky130_fd_sc_hd__nor2_4
X_20529_ _20529_/A _23921_/Q VGND VGND VPWR VPWR _20529_/X sky130_fd_sc_hd__and2_4
XFILLER_126_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24297_ _25526_/CLK _17638_/X HRESETn VGND VGND VPWR VPWR _24297_/Q sky130_fd_sc_hd__dfrtp_4
X_14050_ _14041_/Y _14043_/Y _14046_/Y _14049_/X VGND VGND VPWR VPWR _14050_/X sky130_fd_sc_hd__or4_4
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23248_ _24732_/Q _21021_/X _21024_/X _23247_/X VGND VGND VPWR VPWR _23248_/X sky130_fd_sc_hd__a211o_4
XFILLER_88_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13001_ _13012_/A _13023_/A _13001_/C _13001_/D VGND VGND VPWR VPWR _13001_/X sky130_fd_sc_hd__or4_4
XANTENNA__18446__A1_N _16189_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24419__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23179_ _23095_/X _23178_/X _23141_/X _24834_/Q _23097_/X VGND VGND VPWR VPWR _23180_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_45_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17740_ _17740_/A VGND VGND VPWR VPWR _17762_/A sky130_fd_sc_hd__inv_2
X_14952_ _15241_/A VGND VGND VPWR VPWR _15068_/A sky130_fd_sc_hd__inv_2
XANTENNA__24072__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13903_ _13909_/C VGND VGND VPWR VPWR _13905_/C sky130_fd_sc_hd__buf_2
XANTENNA__18251__B1 _17424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17671_ _17574_/Y _17673_/B _17670_/Y VGND VGND VPWR VPWR _17671_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24001__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14883_ _14882_/X VGND VGND VPWR VPWR _14883_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16278__A _24630_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19410_ _23737_/Q VGND VGND VPWR VPWR _19410_/Y sky130_fd_sc_hd__inv_2
X_16622_ _16622_/A VGND VGND VPWR VPWR _16622_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13834_ _13575_/Y _13829_/X _11829_/X _13833_/X VGND VGND VPWR VPWR _13834_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19341_ _18083_/B VGND VGND VPWR VPWR _19341_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14713__A1_N _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21689__A1 _21682_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13765_ _13748_/C VGND VGND VPWR VPWR _20043_/C sky130_fd_sc_hd__buf_2
X_16553_ _24530_/Q VGND VGND VPWR VPWR _16553_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25278__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18493__A _18414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17010__A1_N _24725_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15504_ _15490_/X VGND VGND VPWR VPWR _15504_/X sky130_fd_sc_hd__buf_2
XANTENNA__22727__B _22727_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12716_ _12707_/A _12707_/B VGND VGND VPWR VPWR _12716_/Y sky130_fd_sc_hd__nand2_4
X_19272_ _19270_/Y _19266_/X _16872_/X _19271_/X VGND VGND VPWR VPWR _23786_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13696_ _13695_/X VGND VGND VPWR VPWR _13696_/Y sky130_fd_sc_hd__inv_2
X_16484_ _16483_/Y _16479_/X _16398_/X _16479_/X VGND VGND VPWR VPWR _16484_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15907__A3 _15768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16725__B _16725_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18223_ _18191_/A _18223_/B _18222_/X VGND VGND VPWR VPWR _18223_/X sky130_fd_sc_hd__and3_4
X_12647_ _12620_/X _12629_/X _12524_/Y VGND VGND VPWR VPWR _12647_/X sky130_fd_sc_hd__o21a_4
X_15435_ _15435_/A _15434_/X VGND VGND VPWR VPWR _15435_/X sky130_fd_sc_hd__or2_4
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15366_ _15369_/A _15369_/B VGND VGND VPWR VPWR _15370_/B sky130_fd_sc_hd__or2_4
X_18154_ _18186_/A _23831_/Q VGND VGND VPWR VPWR _18154_/X sky130_fd_sc_hd__or2_4
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16317__B1 _15959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12578_ _12578_/A _12573_/X _12575_/X _12578_/D VGND VGND VPWR VPWR _12599_/B sky130_fd_sc_hd__or4_4
XFILLER_106_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17105_ _17105_/A _17105_/B VGND VGND VPWR VPWR _17105_/X sky130_fd_sc_hd__or2_4
X_14317_ _25161_/Q _14299_/Y _25160_/Q _14296_/B VGND VGND VPWR VPWR _14317_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17837__A _17837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15297_ _15367_/A _15369_/A _15296_/X VGND VGND VPWR VPWR _15298_/C sky130_fd_sc_hd__or3_4
X_18085_ _18005_/A _18083_/X _18085_/C VGND VGND VPWR VPWR _18086_/C sky130_fd_sc_hd__and3_4
XFILLER_89_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22462__B _22462_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14248_ _13970_/A _13949_/X _13960_/Y _13964_/B VGND VGND VPWR VPWR _14248_/X sky130_fd_sc_hd__or4_4
X_17036_ _17036_/A VGND VGND VPWR VPWR _17036_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24842__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14179_ _14177_/Y _14110_/X _14136_/X _14178_/Y VGND VGND VPWR VPWR _14179_/X sky130_fd_sc_hd__o22a_4
XFILLER_97_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18987_ _19152_/A _14671_/X _25061_/Q _18987_/D VGND VGND VPWR VPWR _18987_/X sky130_fd_sc_hd__or4_4
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17938_ _17956_/A _23828_/Q VGND VGND VPWR VPWR _17939_/C sky130_fd_sc_hd__or2_4
XFILLER_85_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17869_ _16911_/Y _17867_/X _17868_/Y VGND VGND VPWR VPWR _24252_/D sky130_fd_sc_hd__o21a_4
XANTENNA__18793__A1 _18608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19608_ _23668_/Q VGND VGND VPWR VPWR _19608_/Y sky130_fd_sc_hd__inv_2
X_20880_ _20877_/Y _20878_/Y _20879_/X VGND VGND VPWR VPWR _20880_/X sky130_fd_sc_hd__o21a_4
X_19539_ _19538_/X VGND VGND VPWR VPWR _19539_/X sky130_fd_sc_hd__buf_2
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22550_ _22550_/A _22590_/B VGND VGND VPWR VPWR _22550_/X sky130_fd_sc_hd__or2_4
XFILLER_62_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16556__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18860__A2_N _18789_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21501_ _21162_/X VGND VGND VPWR VPWR _21502_/A sky130_fd_sc_hd__buf_2
X_22481_ _22476_/X _22478_/X _22479_/X _24712_/Q _22480_/X VGND VGND VPWR VPWR _22482_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24220_ _24219_/CLK _18248_/X HRESETn VGND VGND VPWR VPWR _24220_/Q sky130_fd_sc_hd__dfrtp_4
X_21432_ _21293_/A VGND VGND VPWR VPWR _22590_/B sky130_fd_sc_hd__buf_2
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12593__B2 _24872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24151_ _24151_/CLK _24151_/D HRESETn VGND VGND VPWR VPWR _18393_/A sky130_fd_sc_hd__dfrtp_4
X_21363_ _23670_/Q _21362_/X _19555_/Y _21362_/X VGND VGND VPWR VPWR _21363_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17747__A _17744_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23102_ _21418_/X VGND VGND VPWR VPWR _23102_/X sky130_fd_sc_hd__buf_2
X_20314_ _20313_/Y _20311_/X _19995_/X _20311_/X VGND VGND VPWR VPWR _20314_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21269__A _13593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24082_ _24398_/CLK _20952_/X HRESETn VGND VGND VPWR VPWR RsTx_S0 sky130_fd_sc_hd__dfstp_4
X_21294_ _24600_/Q _21293_/X VGND VGND VPWR VPWR _21294_/X sky130_fd_sc_hd__or2_4
XANTENNA__24583__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23033_ _23143_/A _23033_/B VGND VGND VPWR VPWR _23033_/X sky130_fd_sc_hd__and2_4
X_20245_ _20232_/Y VGND VGND VPWR VPWR _20245_/X sky130_fd_sc_hd__buf_2
XFILLER_116_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24512__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20176_ _20174_/Y _20170_/X _20085_/X _20175_/X VGND VGND VPWR VPWR _23466_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24984_ _24984_/CLK _15357_/X HRESETn VGND VGND VPWR VPWR _24984_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23935_ _25122_/CLK _23935_/D HRESETn VGND VGND VPWR VPWR _18873_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22580__A2 _22534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13515__A _11862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11880_ _11700_/X VGND VGND VPWR VPWR _11880_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23866_ _25485_/CLK _19046_/X VGND VGND VPWR VPWR _19044_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__25371__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22817_ _24720_/Q _21049_/X _21050_/X _22816_/X VGND VGND VPWR VPWR _22817_/X sky130_fd_sc_hd__a211o_4
XFILLER_60_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23797_ _23798_/CLK _19240_/X VGND VGND VPWR VPWR _13436_/B sky130_fd_sc_hd__dfxtp_4
X_13550_ _13551_/A _14598_/A _13549_/Y _13582_/A VGND VGND VPWR VPWR _13550_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25300__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25536_ _24691_/CLK _25536_/D HRESETn VGND VGND VPWR VPWR _25536_/Q sky130_fd_sc_hd__dfrtp_4
X_22748_ _16682_/Y _22598_/B VGND VGND VPWR VPWR _22748_/X sky130_fd_sc_hd__and2_4
X_12501_ _12264_/X _12499_/X _12500_/Y VGND VGND VPWR VPWR _12501_/X sky130_fd_sc_hd__o21a_4
X_13481_ _13481_/A VGND VGND VPWR VPWR _13481_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25467_ _24097_/CLK _25467_/D HRESETn VGND VGND VPWR VPWR _12088_/A sky130_fd_sc_hd__dfrtp_4
X_22679_ _22782_/A _22679_/B VGND VGND VPWR VPWR _22679_/Y sky130_fd_sc_hd__nor2_4
X_15220_ _14926_/X _15219_/X _15174_/X VGND VGND VPWR VPWR _15220_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_55_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12432_ _12432_/A _12432_/B VGND VGND VPWR VPWR _12433_/B sky130_fd_sc_hd__or2_4
X_24418_ _24431_/CLK _16822_/X HRESETn VGND VGND VPWR VPWR _24418_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23293__B1 _22834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18839__A2 _18630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25398_ _25411_/CLK _25398_/D HRESETn VGND VGND VPWR VPWR _25398_/Q sky130_fd_sc_hd__dfrtp_4
X_15151_ _24985_/Q _15149_/Y _15298_/B _15147_/A VGND VGND VPWR VPWR _15152_/D sky130_fd_sc_hd__a2bb2o_4
X_12363_ _25326_/Q VGND VGND VPWR VPWR _12363_/Y sky130_fd_sc_hd__inv_2
X_24349_ _24345_/CLK _24349_/D HRESETn VGND VGND VPWR VPWR _17177_/A sky130_fd_sc_hd__dfrtp_4
X_14102_ _14102_/A _14102_/B _14117_/A VGND VGND VPWR VPWR _14103_/B sky130_fd_sc_hd__or3_4
X_15082_ _15074_/X _15082_/B _15079_/X _15082_/D VGND VGND VPWR VPWR _15121_/A sky130_fd_sc_hd__or4_4
XANTENNA__23045__B1 _25530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12294_ _25353_/Q VGND VGND VPWR VPWR _12294_/Y sky130_fd_sc_hd__inv_2
X_14033_ _14042_/A _14003_/C VGND VGND VPWR VPWR _14045_/A sky130_fd_sc_hd__or2_4
X_18910_ _18909_/Y _18907_/X _16876_/X _18907_/X VGND VGND VPWR VPWR _23913_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22399__A2 _18272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19890_ _19902_/A VGND VGND VPWR VPWR _19890_/X sky130_fd_sc_hd__buf_2
XANTENNA__24253__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18841_ _24564_/Q _18671_/A _16463_/Y _18698_/C VGND VGND VPWR VPWR _18843_/C sky130_fd_sc_hd__o22a_4
XFILLER_136_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18772_ _18772_/A _18693_/A VGND VGND VPWR VPWR _18773_/B sky130_fd_sc_hd__or2_4
XFILLER_121_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15984_ _15788_/X _15857_/A _15836_/X _24739_/Q _15933_/A VGND VGND VPWR VPWR _15984_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_94_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17723_ _24205_/Q _17710_/X VGND VGND VPWR VPWR _17724_/A sky130_fd_sc_hd__and2_4
X_14935_ _25004_/Q _14934_/A _15262_/A _14934_/Y VGND VGND VPWR VPWR _14939_/C sky130_fd_sc_hd__o22a_4
XFILLER_110_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25459__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13425__A _13457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17654_ _17571_/Y _17653_/X VGND VGND VPWR VPWR _17657_/B sky130_fd_sc_hd__or2_4
X_14866_ _14865_/X VGND VGND VPWR VPWR _14866_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16605_ _16603_/Y _16601_/X _16604_/X _16601_/X VGND VGND VPWR VPWR _24510_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13817_ _13817_/A VGND VGND VPWR VPWR _21994_/A sky130_fd_sc_hd__buf_2
X_17585_ _17585_/A _17585_/B VGND VGND VPWR VPWR _17586_/B sky130_fd_sc_hd__nor2_4
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14797_ _25042_/Q VGND VGND VPWR VPWR _14819_/C sky130_fd_sc_hd__inv_2
XFILLER_17_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19324_ _23767_/Q VGND VGND VPWR VPWR _19324_/Y sky130_fd_sc_hd__inv_2
X_16536_ _16535_/Y _16531_/X _16442_/X _16531_/X VGND VGND VPWR VPWR _24536_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19112__A _19106_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25041__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13748_ _13748_/A _13763_/A _13748_/C _13754_/A VGND VGND VPWR VPWR _13748_/X sky130_fd_sc_hd__and4_4
XANTENNA__16538__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16455__B _16725_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19255_ _19255_/A VGND VGND VPWR VPWR _21598_/B sky130_fd_sc_hd__inv_2
XFILLER_108_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16467_ _16474_/A VGND VGND VPWR VPWR _16467_/X sky130_fd_sc_hd__buf_2
X_13679_ _13694_/B VGND VGND VPWR VPWR _13721_/A sky130_fd_sc_hd__inv_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14256__A _21139_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18206_ _17973_/X _18206_/B VGND VGND VPWR VPWR _18208_/B sky130_fd_sc_hd__or2_4
X_15418_ _15416_/Y _15417_/X _15407_/X VGND VGND VPWR VPWR _24966_/D sky130_fd_sc_hd__and3_4
X_19186_ _19185_/Y _19181_/X _19117_/X _19181_/X VGND VGND VPWR VPWR _19186_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_23_0_HCLK clkbuf_5_22_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16398_ HWDATA[22] VGND VGND VPWR VPWR _16398_/X sky130_fd_sc_hd__buf_2
X_18137_ _18137_/A _18135_/X _18136_/X VGND VGND VPWR VPWR _18138_/C sky130_fd_sc_hd__and3_4
XANTENNA__21834__A1 _21106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15349_ _15349_/A VGND VGND VPWR VPWR _24985_/D sky130_fd_sc_hd__inv_2
XFILLER_129_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16471__A _24561_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18068_ _18137_/A _18068_/B _18068_/C VGND VGND VPWR VPWR _18069_/C sky130_fd_sc_hd__and3_4
XFILLER_117_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16710__B1 _16355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14703__B _14675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17019_ _17346_/B VGND VGND VPWR VPWR _17260_/A sky130_fd_sc_hd__buf_2
XANTENNA__12504__A _12280_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20030_ _22010_/B _20024_/X _19981_/X _20029_/X VGND VGND VPWR VPWR _23522_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_147_0_HCLK clkbuf_7_73_0_HCLK/X VGND VGND VPWR VPWR _25508_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__23976__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21981_ _22035_/A _21980_/X _21502_/X VGND VGND VPWR VPWR _21981_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_66_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23720_ _23887_/CLK _19457_/X VGND VGND VPWR VPWR _18110_/B sky130_fd_sc_hd__dfxtp_4
X_20932_ _20929_/Y _20930_/Y _20931_/X VGND VGND VPWR VPWR _20932_/X sky130_fd_sc_hd__o21a_4
XFILLER_54_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16777__B1 _16521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23651_ _23649_/CLK _19667_/X VGND VGND VPWR VPWR _23651_/Q sky130_fd_sc_hd__dfxtp_4
X_20863_ _20863_/A VGND VGND VPWR VPWR _20913_/A sky130_fd_sc_hd__inv_2
XFILLER_74_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22602_ _22602_/A VGND VGND VPWR VPWR _22602_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16529__B1 _16528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23582_ _24089_/CLK _23582_/D VGND VGND VPWR VPWR _23582_/Q sky130_fd_sc_hd__dfxtp_4
X_20794_ _20770_/X _20793_/X _15572_/A _20774_/X VGND VGND VPWR VPWR _24023_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25321_ _24840_/CLK _25321_/D HRESETn VGND VGND VPWR VPWR _21007_/A sky130_fd_sc_hd__dfrtp_4
X_22533_ _21270_/X _22531_/X _21950_/X _22532_/X VGND VGND VPWR VPWR _22533_/X sky130_fd_sc_hd__o22a_4
X_25252_ _25279_/CLK _13830_/X HRESETn VGND VGND VPWR VPWR _13580_/A sky130_fd_sc_hd__dfrtp_4
X_22464_ _22464_/A VGND VGND VPWR VPWR _23304_/B sky130_fd_sc_hd__buf_2
XANTENNA__24764__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24203_ _24288_/CLK _24203_/D HRESETn VGND VGND VPWR VPWR _17713_/A sky130_fd_sc_hd__dfrtp_4
X_21415_ _21284_/A VGND VGND VPWR VPWR _21416_/A sky130_fd_sc_hd__buf_2
XANTENNA__12566__B2 _24854_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21825__B2 _22873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25183_ _25192_/CLK _14237_/X HRESETn VGND VGND VPWR VPWR _25183_/Q sky130_fd_sc_hd__dfstp_4
X_22395_ _22395_/A _21026_/B VGND VGND VPWR VPWR _22395_/X sky130_fd_sc_hd__or2_4
XFILLER_120_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24134_ _24133_/CLK _24134_/D HRESETn VGND VGND VPWR VPWR _18610_/A sky130_fd_sc_hd__dfrtp_4
X_21346_ _18386_/Y _16453_/B _12166_/A _12096_/X VGND VGND VPWR VPWR _21346_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16701__B1 _16604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24065_ _24715_/CLK _20461_/X HRESETn VGND VGND VPWR VPWR _24065_/Q sky130_fd_sc_hd__dfrtp_4
X_21277_ _22827_/A VGND VGND VPWR VPWR _21277_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12414__A _12252_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23016_ _21409_/A _23014_/Y _22826_/X _23015_/X VGND VGND VPWR VPWR _23017_/A sky130_fd_sc_hd__o22a_4
X_20228_ _23445_/Q VGND VGND VPWR VPWR _20228_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_43_0_HCLK clkbuf_7_42_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_87_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15268__B1 _15174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15725__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20159_ _20158_/Y _20154_/X _20092_/X _20154_/X VGND VGND VPWR VPWR _23472_/D sky130_fd_sc_hd__a2bb2o_4
X_12981_ _21006_/A _12866_/X _12980_/Y VGND VGND VPWR VPWR _25354_/D sky130_fd_sc_hd__o21a_4
XFILLER_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24967_ _24977_/CLK _15413_/Y HRESETn VGND VGND VPWR VPWR _15144_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23315__A1_N _17264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14720_ _14719_/X VGND VGND VPWR VPWR _14720_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13245__A _13156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11932_ _11932_/A VGND VGND VPWR VPWR _19618_/A sky130_fd_sc_hd__buf_2
X_23918_ _23978_/CLK _20967_/X HRESETn VGND VGND VPWR VPWR _22097_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16768__B1 _15750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24898_ _24868_/CLK _15594_/X HRESETn VGND VGND VPWR VPWR _24898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_72_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11863_ _11860_/Y _11741_/X _11862_/X _11741_/X VGND VGND VPWR VPWR _11863_/X sky130_fd_sc_hd__a2bb2o_4
X_14651_ _18010_/A VGND VGND VPWR VPWR _17930_/A sky130_fd_sc_hd__buf_2
X_23849_ _24396_/CLK _23849_/D VGND VGND VPWR VPWR _23849_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13602_ _13624_/A VGND VGND VPWR VPWR _18987_/D sky130_fd_sc_hd__buf_2
X_17370_ _17370_/A _17370_/B _17369_/Y VGND VGND VPWR VPWR _17370_/X sky130_fd_sc_hd__and3_4
XFILLER_60_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11794_ _11750_/A VGND VGND VPWR VPWR _11794_/X sky130_fd_sc_hd__buf_2
X_14582_ _13568_/X _14582_/B VGND VGND VPWR VPWR _14582_/X sky130_fd_sc_hd__or2_4
XFILLER_92_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20316__B2 _20298_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20078__A _20095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16321_ _16320_/Y _16316_/X _15964_/X _16316_/X VGND VGND VPWR VPWR _24616_/D sky130_fd_sc_hd__a2bb2o_4
X_13533_ _13533_/A _13533_/B _15652_/D _13533_/D VGND VGND VPWR VPWR _13534_/A sky130_fd_sc_hd__or4_4
X_25519_ _24275_/CLK _11814_/X HRESETn VGND VGND VPWR VPWR _25519_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19040_ _19052_/A VGND VGND VPWR VPWR _19040_/X sky130_fd_sc_hd__buf_2
X_13464_ _13196_/Y _13463_/X _25313_/Q _13195_/X VGND VGND VPWR VPWR _13464_/X sky130_fd_sc_hd__o22a_4
X_16252_ _16251_/Y _16247_/X _16057_/X _16247_/X VGND VGND VPWR VPWR _16252_/X sky130_fd_sc_hd__a2bb2o_4
X_12415_ _12244_/Y _12414_/X VGND VGND VPWR VPWR _12415_/X sky130_fd_sc_hd__or2_4
X_15203_ _25018_/Q _15203_/B VGND VGND VPWR VPWR _15203_/X sky130_fd_sc_hd__or2_4
XFILLER_127_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17387__A _17387_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13395_ _13395_/A _23599_/Q VGND VGND VPWR VPWR _13395_/X sky130_fd_sc_hd__or2_4
X_16183_ _16183_/A _22444_/A VGND VGND VPWR VPWR _16184_/A sky130_fd_sc_hd__or2_4
XANTENNA__24434__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12346_ _25323_/Q _12344_/Y _13102_/A _12345_/Y VGND VGND VPWR VPWR _12346_/X sky130_fd_sc_hd__a2bb2o_4
X_15134_ _15133_/Y _16421_/A _15133_/Y _16421_/A VGND VGND VPWR VPWR _15134_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15950__A1_N _12207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13506__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15065_ _15065_/A VGND VGND VPWR VPWR _15065_/Y sky130_fd_sc_hd__inv_2
X_19942_ _19942_/A VGND VGND VPWR VPWR _19942_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12277_ _12277_/A _12277_/B VGND VGND VPWR VPWR _12289_/C sky130_fd_sc_hd__or2_4
XANTENNA__12324__A _24814_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22740__B _22626_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14016_ _25216_/Q _13985_/B VGND VGND VPWR VPWR _14016_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__18445__B1 _21322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19873_ _19880_/A VGND VGND VPWR VPWR _19873_/X sky130_fd_sc_hd__buf_2
XFILLER_122_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18824_ _16493_/Y _24131_/Q _16493_/Y _24131_/Q VGND VGND VPWR VPWR _18828_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19107__A _19106_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15965__A1_N _12228_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12978__B _12631_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18755_ _18626_/Y _18759_/B _18754_/Y VGND VGND VPWR VPWR _24132_/D sky130_fd_sc_hd__o21a_4
XANTENNA__14896__D _14895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25293__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_0_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15967_ _15967_/A VGND VGND VPWR VPWR _15967_/X sky130_fd_sc_hd__buf_2
XFILLER_76_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18946__A _18945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17706_ _17706_/A VGND VGND VPWR VPWR _21467_/A sky130_fd_sc_hd__buf_2
XFILLER_48_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14918_ _25019_/Q VGND VGND VPWR VPWR _15194_/A sky130_fd_sc_hd__inv_2
XANTENNA__25222__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18686_ _18686_/A VGND VGND VPWR VPWR _18692_/B sky130_fd_sc_hd__inv_2
X_15898_ _12755_/Y _15896_/X _15897_/X _15896_/X VGND VGND VPWR VPWR _24782_/D sky130_fd_sc_hd__a2bb2o_4
X_17637_ _17567_/A _17642_/B _17590_/X VGND VGND VPWR VPWR _17637_/Y sky130_fd_sc_hd__a21oi_4
X_14849_ _14815_/C _14801_/B _14815_/C _14801_/B VGND VGND VPWR VPWR _14849_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22187__B _22157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12245__B1 _12244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17568_ _17521_/Y _17525_/Y _17567_/X VGND VGND VPWR VPWR _17568_/X sky130_fd_sc_hd__or3_4
X_19307_ _17442_/X VGND VGND VPWR VPWR _19307_/X sky130_fd_sc_hd__buf_2
X_16519_ _16518_/Y _16516_/X _16147_/X _16516_/X VGND VGND VPWR VPWR _24542_/D sky130_fd_sc_hd__a2bb2o_4
X_17499_ _24288_/Q VGND VGND VPWR VPWR _17499_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19238_ _19237_/Y _19235_/X _19191_/X _19235_/X VGND VGND VPWR VPWR _19238_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16931__B1 _16130_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18830__A1_N _16539_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19169_ _19169_/A VGND VGND VPWR VPWR _19169_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21200_ _21200_/A _21200_/B VGND VGND VPWR VPWR _21200_/X sky130_fd_sc_hd__or2_4
XANTENNA__16540__A2_N _16461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22180_ _21043_/Y VGND VGND VPWR VPWR _22186_/A sky130_fd_sc_hd__buf_2
XANTENNA__24104__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21131_ _25475_/Q _13789_/B _23343_/B _12059_/X VGND VGND VPWR VPWR _21131_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18845__A1_N _24539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21062_ _15784_/B VGND VGND VPWR VPWR _21062_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20243__B1 _19740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20013_ _20013_/A VGND VGND VPWR VPWR _20013_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19017__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20794__B2 _20774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24821_ _24821_/CLK _15821_/X HRESETn VGND VGND VPWR VPWR _24821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17760__A _17751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21964_ _21960_/Y _21961_/X _21962_/X _21963_/X VGND VGND VPWR VPWR _21964_/X sky130_fd_sc_hd__a211o_4
XFILLER_27_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24752_ _24759_/CLK _15965_/X HRESETn VGND VGND VPWR VPWR _24752_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21743__B1 _21587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20915_ _20889_/B _13650_/X VGND VGND VPWR VPWR _20915_/Y sky130_fd_sc_hd__nor2_4
X_23703_ _23398_/CLK _19508_/X VGND VGND VPWR VPWR _19506_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_27_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24683_ _24682_/CLK _16129_/X HRESETn VGND VGND VPWR VPWR _22745_/A sky130_fd_sc_hd__dfrtp_4
X_21895_ _21614_/A _21884_/X _21894_/X VGND VGND VPWR VPWR _21895_/X sky130_fd_sc_hd__or3_4
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16376__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22299__A1 _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23634_ _23649_/CLK _19713_/X VGND VGND VPWR VPWR _23634_/Q sky130_fd_sc_hd__dfxtp_4
X_20846_ _13659_/A VGND VGND VPWR VPWR _20846_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23565_ _24309_/CLK _23565_/D VGND VGND VPWR VPWR _19906_/A sky130_fd_sc_hd__dfxtp_4
X_20777_ _24019_/Q _20772_/X _20776_/Y VGND VGND VPWR VPWR _20777_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_70_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22516_ _22515_/X VGND VGND VPWR VPWR _22782_/A sky130_fd_sc_hd__buf_2
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25304_ _25305_/CLK _25304_/D HRESETn VGND VGND VPWR VPWR _25304_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23248__B1 _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23496_ _23496_/CLK _23496_/D VGND VGND VPWR VPWR _23496_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22447_ _15668_/X _22447_/B VGND VGND VPWR VPWR _22447_/Y sky130_fd_sc_hd__nor2_4
XFILLER_10_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25235_ _25172_/CLK _13875_/X HRESETn VGND VGND VPWR VPWR _21829_/A sky130_fd_sc_hd__dfrtp_4
X_12200_ _22853_/A VGND VGND VPWR VPWR _12200_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23263__A3 _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13180_ _13180_/A _13180_/B VGND VGND VPWR VPWR _13180_/X sky130_fd_sc_hd__or2_4
XFILLER_100_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25166_ _25305_/CLK _14304_/Y HRESETn VGND VGND VPWR VPWR _12027_/D sky130_fd_sc_hd__dfrtp_4
X_22378_ _21890_/X _22374_/X _22375_/X _22376_/X _22377_/X VGND VGND VPWR VPWR _22378_/X
+ sky130_fd_sc_hd__a32o_4
X_12131_ _12106_/Y _12130_/X VGND VGND VPWR VPWR _12131_/Y sky130_fd_sc_hd__nor2_4
XFILLER_123_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20482__B1 _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24117_ _24117_/CLK _18812_/Y HRESETn VGND VGND VPWR VPWR _24117_/Q sky130_fd_sc_hd__dfrtp_4
X_21329_ _16451_/A _21322_/X _21329_/C VGND VGND VPWR VPWR _21407_/B sky130_fd_sc_hd__and3_4
XFILLER_2_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25097_ _24077_/CLK _25097_/D HRESETn VGND VGND VPWR VPWR _20441_/B sky130_fd_sc_hd__dfrtp_4
X_12062_ _12046_/Y _12061_/Y _11867_/X _12061_/Y VGND VGND VPWR VPWR _12062_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14161__B1 _25122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24048_ _24049_/CLK _20904_/Y HRESETn VGND VGND VPWR VPWR _13649_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_104_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20234__B1 _18247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16870_ _20089_/A VGND VGND VPWR VPWR _19787_/A sky130_fd_sc_hd__buf_2
XFILLER_133_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20785__B2 _20774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15821_ _15816_/X _15819_/X _15745_/X _24821_/Q _15817_/X VGND VGND VPWR VPWR _15821_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_130_0_HCLK clkbuf_7_65_0_HCLK/X VGND VGND VPWR VPWR _23446_/CLK sky130_fd_sc_hd__clkbuf_1
X_18540_ _18540_/A _18540_/B VGND VGND VPWR VPWR _18540_/Y sky130_fd_sc_hd__nand2_4
X_15752_ HWDATA[11] VGND VGND VPWR VPWR _15752_/X sky130_fd_sc_hd__buf_2
X_12964_ _12964_/A _12964_/B _12963_/Y VGND VGND VPWR VPWR _25361_/D sky130_fd_sc_hd__and3_4
Xclkbuf_8_193_0_HCLK clkbuf_7_96_0_HCLK/X VGND VGND VPWR VPWR _24177_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14703_ _14703_/A _14675_/X _14698_/X _14702_/X VGND VGND VPWR VPWR _14703_/X sky130_fd_sc_hd__or4_4
XANTENNA__21192__A _21192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11915_ _11877_/A _11914_/X _11912_/Y VGND VGND VPWR VPWR _11915_/X sky130_fd_sc_hd__o21a_4
X_18471_ _24156_/Q VGND VGND VPWR VPWR _18471_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22719__C _22711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15683_ _15682_/X VGND VGND VPWR VPWR _15683_/Y sky130_fd_sc_hd__inv_2
X_12895_ _12886_/X VGND VGND VPWR VPWR _12896_/B sky130_fd_sc_hd__inv_2
X_17422_ _17420_/Y _17417_/X _17421_/X _17417_/X VGND VGND VPWR VPWR _24319_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15190__A _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14634_ _14632_/A VGND VGND VPWR VPWR _14634_/Y sky130_fd_sc_hd__inv_2
X_11846_ _15766_/A VGND VGND VPWR VPWR _16355_/A sky130_fd_sc_hd__buf_2
XANTENNA__24686__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17353_ _17240_/Y _17353_/B VGND VGND VPWR VPWR _17354_/C sky130_fd_sc_hd__or2_4
XANTENNA__21920__A _21942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11777_ _11777_/A VGND VGND VPWR VPWR _11777_/X sky130_fd_sc_hd__buf_2
X_14565_ _14598_/A _14564_/X VGND VGND VPWR VPWR _14596_/B sky130_fd_sc_hd__or2_4
XANTENNA__24615__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16304_ _16302_/Y _16296_/X _15949_/X _16303_/X VGND VGND VPWR VPWR _24623_/D sky130_fd_sc_hd__a2bb2o_4
X_13516_ _13514_/Y _13512_/X _13515_/X _13512_/X VGND VGND VPWR VPWR _25295_/D sky130_fd_sc_hd__a2bb2o_4
X_17284_ _24355_/Q _17284_/B VGND VGND VPWR VPWR _17286_/B sky130_fd_sc_hd__or2_4
X_14496_ _14036_/A _23922_/Q VGND VGND VPWR VPWR _14496_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_4_1_0_HCLK_A clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19023_ _19030_/A VGND VGND VPWR VPWR _19023_/X sky130_fd_sc_hd__buf_2
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16235_ _11809_/A VGND VGND VPWR VPWR _16235_/X sky130_fd_sc_hd__buf_2
X_13447_ _13297_/X _13439_/X _13447_/C VGND VGND VPWR VPWR _13447_/X sky130_fd_sc_hd__and3_4
XANTENNA__20068__A3 _11838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13378_ _13309_/A _13378_/B _13377_/X VGND VGND VPWR VPWR _13378_/X sky130_fd_sc_hd__and3_4
X_16166_ _16165_/Y _16088_/A _15480_/X _16088_/A VGND VGND VPWR VPWR _24668_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13795__D _13795_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18130__A2 _18114_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12950__A1 _12944_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15117_ _24981_/Q VGND VGND VPWR VPWR _15367_/A sky130_fd_sc_hd__inv_2
X_12329_ _25351_/Q _24836_/Q _13001_/C _12328_/Y VGND VGND VPWR VPWR _12339_/A sky130_fd_sc_hd__o22a_4
X_16097_ _16096_/Y _16094_/X _15942_/X _16094_/X VGND VGND VPWR VPWR _16097_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12054__A _12054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15048_ _14886_/X _24444_/Q _14966_/A _15027_/Y VGND VGND VPWR VPWR _15054_/A sky130_fd_sc_hd__a2bb2o_4
X_19925_ _19925_/A VGND VGND VPWR VPWR _19925_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25474__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20225__B1 _19721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19856_ _23584_/Q VGND VGND VPWR VPWR _21764_/B sky130_fd_sc_hd__inv_2
XANTENNA__25403__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18807_ _18799_/A _18803_/X _18806_/Y VGND VGND VPWR VPWR _18807_/X sky130_fd_sc_hd__and3_4
XFILLER_56_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19787_ _19787_/A VGND VGND VPWR VPWR _19787_/X sky130_fd_sc_hd__buf_2
X_16999_ _16042_/Y _17036_/A _16042_/Y _17036_/A VGND VGND VPWR VPWR _17003_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18738_ _18738_/A _18728_/B _18738_/C VGND VGND VPWR VPWR _18738_/X sky130_fd_sc_hd__and3_4
X_18669_ _18669_/A VGND VGND VPWR VPWR _18742_/A sky130_fd_sc_hd__buf_2
XFILLER_110_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20700_ _20699_/Y _20694_/Y _13128_/B VGND VGND VPWR VPWR _20700_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12218__B1 _12385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21680_ _21675_/X _21678_/X _21679_/X VGND VGND VPWR VPWR _21681_/C sky130_fd_sc_hd__o21a_4
X_20631_ _15461_/Y _20628_/X _20619_/X _20630_/X VGND VGND VPWR VPWR _20632_/A sky130_fd_sc_hd__a211o_4
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24356__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23350_ VGND VGND VPWR VPWR _23350_/HI scl_o_S4 sky130_fd_sc_hd__conb_1
X_20562_ _20562_/A VGND VGND VPWR VPWR _20571_/C sky130_fd_sc_hd__buf_2
XFILLER_137_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22301_ _23170_/A _22301_/B _22301_/C VGND VGND VPWR VPWR _22301_/X sky130_fd_sc_hd__and3_4
X_23281_ _23281_/A _23281_/B _23281_/C _23280_/X VGND VGND VPWR VPWR _23281_/X sky130_fd_sc_hd__or4_4
X_20493_ _20493_/A _20602_/A _20479_/C VGND VGND VPWR VPWR _20493_/X sky130_fd_sc_hd__and3_4
XANTENNA__14444__A _25121_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25020_ _25020_/CLK _15198_/X HRESETn VGND VGND VPWR VPWR _25020_/Q sky130_fd_sc_hd__dfrtp_4
X_22232_ _22247_/A _22229_/X _22231_/X VGND VGND VPWR VPWR _22232_/X sky130_fd_sc_hd__and3_4
XANTENNA__22453__A1 _22613_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18657__B1 _24522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22453__B2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22163_ _22162_/X VGND VGND VPWR VPWR _22163_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23991__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21114_ _21408_/A _21108_/X _21114_/C VGND VGND VPWR VPWR _21114_/X sky130_fd_sc_hd__and3_4
XFILLER_117_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22094_ _20452_/A _21843_/X VGND VGND VPWR VPWR _22101_/A sky130_fd_sc_hd__nor2_4
XFILLER_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23920__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15891__B1 _22708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21045_ _22146_/A VGND VGND VPWR VPWR _21045_/X sky130_fd_sc_hd__buf_2
XANTENNA__25144__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24804_ _24804_/CLK _24804_/D HRESETn VGND VGND VPWR VPWR _12980_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_203_0_HCLK clkbuf_8_203_0_HCLK/A VGND VGND VPWR VPWR _24804_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22996_ _15089_/A _23171_/B VGND VGND VPWR VPWR _23001_/B sky130_fd_sc_hd__or2_4
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_9_0_HCLK clkbuf_7_4_0_HCLK/X VGND VGND VPWR VPWR _23467_/CLK sky130_fd_sc_hd__clkbuf_1
X_24735_ _24811_/CLK _24735_/D HRESETn VGND VGND VPWR VPWR _24735_/Q sky130_fd_sc_hd__dfrtp_4
X_21947_ _21943_/X _21946_/X _18298_/X VGND VGND VPWR VPWR _21948_/C sky130_fd_sc_hd__o21a_4
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11666_/X _11700_/B _11688_/X _11699_/X VGND VGND VPWR VPWR _11700_/X sky130_fd_sc_hd__or4_4
XFILLER_128_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12683_/A _12686_/B VGND VGND VPWR VPWR _12684_/B sky130_fd_sc_hd__or2_4
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ _21904_/A _19251_/Y VGND VGND VPWR VPWR _21878_/X sky130_fd_sc_hd__or2_4
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24666_ _23467_/CLK _24666_/D HRESETn VGND VGND VPWR VPWR _13744_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _20828_/Y _13654_/A _13656_/B VGND VGND VPWR VPWR _20829_/X sky130_fd_sc_hd__o21a_4
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23617_ _23683_/CLK _19762_/X VGND VGND VPWR VPWR _23617_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24097__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16834__A _24413_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24597_ _24596_/CLK _24597_/D HRESETn VGND VGND VPWR VPWR _16378_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14350_ _24094_/Q _14345_/X _14349_/X VGND VGND VPWR VPWR _14350_/X sky130_fd_sc_hd__and3_4
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18896__B1 _17443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24026__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23548_ _23545_/CLK _23548_/D VGND VGND VPWR VPWR _19949_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13301_ _13155_/Y VGND VGND VPWR VPWR _13301_/X sky130_fd_sc_hd__buf_2
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14281_ _20515_/B VGND VGND VPWR VPWR _14281_/X sky130_fd_sc_hd__buf_2
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23479_ _23478_/CLK _20141_/X VGND VGND VPWR VPWR _20139_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_7_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13232_ _17453_/A VGND VGND VPWR VPWR _13390_/A sky130_fd_sc_hd__buf_2
X_16020_ _16019_/Y _16015_/X _15952_/X _16015_/X VGND VGND VPWR VPWR _16020_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18648__B1 _16565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25218_ _25219_/CLK _14086_/X HRESETn VGND VGND VPWR VPWR _14002_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13163_ _13154_/X _13160_/X _13162_/X VGND VGND VPWR VPWR _13163_/X sky130_fd_sc_hd__o21a_4
X_25149_ _24109_/CLK _14353_/Y HRESETn VGND VGND VPWR VPWR _14339_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_87_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12114_ _12119_/A VGND VGND VPWR VPWR _12114_/X sky130_fd_sc_hd__buf_2
X_13094_ _12991_/B _13097_/B VGND VGND VPWR VPWR _13095_/C sky130_fd_sc_hd__nand2_4
X_17971_ _18087_/A VGND VGND VPWR VPWR _18137_/A sky130_fd_sc_hd__buf_2
XFILLER_97_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17384__B _17384_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19710_ _19709_/Y _19707_/X _19642_/X _19707_/X VGND VGND VPWR VPWR _23635_/D sky130_fd_sc_hd__a2bb2o_4
X_12045_ _24093_/Q _12028_/A _25475_/Q _12041_/X VGND VGND VPWR VPWR _25475_/D sky130_fd_sc_hd__o22a_4
X_16922_ _16922_/A _16922_/B _16922_/C _16922_/D VGND VGND VPWR VPWR _16922_/X sky130_fd_sc_hd__or4_4
XANTENNA__12602__A _12602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_13_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_66_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21955__B1 _23336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19641_ _13242_/B VGND VGND VPWR VPWR _19641_/Y sky130_fd_sc_hd__inv_2
X_16853_ _14937_/Y _16848_/X _16852_/X _16848_/X VGND VGND VPWR VPWR _16853_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21915__A _21942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15804_ _15781_/X _15795_/X _15723_/X _24833_/Q _15793_/X VGND VGND VPWR VPWR _15804_/X
+ sky130_fd_sc_hd__a32o_4
X_19572_ _21810_/B _19567_/X _11948_/X _19567_/X VGND VGND VPWR VPWR _23680_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16784_ _15027_/Y _16778_/X _16782_/X _16783_/X VGND VGND VPWR VPWR _24437_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_24_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13996_ _13990_/C VGND VGND VPWR VPWR _14006_/B sky130_fd_sc_hd__inv_2
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24867__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18523_ _18523_/A _18523_/B VGND VGND VPWR VPWR _18523_/X sky130_fd_sc_hd__or2_4
X_15735_ _15721_/A VGND VGND VPWR VPWR _15735_/X sky130_fd_sc_hd__buf_2
X_12947_ _12842_/A _12945_/A VGND VGND VPWR VPWR _12947_/X sky130_fd_sc_hd__or2_4
XFILLER_59_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18454_ _18521_/A VGND VGND VPWR VPWR _18517_/A sky130_fd_sc_hd__buf_2
XFILLER_45_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15666_ _21556_/A VGND VGND VPWR VPWR _15667_/A sky130_fd_sc_hd__buf_2
X_12878_ _12880_/B VGND VGND VPWR VPWR _12879_/B sky130_fd_sc_hd__inv_2
X_17405_ _17387_/X _17401_/X _24326_/Q _20992_/A _17404_/X VGND VGND VPWR VPWR _17405_/X
+ sky130_fd_sc_hd__a32o_4
X_14617_ _14632_/A _14616_/X VGND VGND VPWR VPWR _14617_/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11829_ HWDATA[8] VGND VGND VPWR VPWR _11829_/X sky130_fd_sc_hd__buf_2
X_18385_ _18383_/Y _18384_/X _24179_/Q _18384_/X VGND VGND VPWR VPWR _24180_/D sky130_fd_sc_hd__a2bb2o_4
X_15597_ _15597_/A VGND VGND VPWR VPWR _22787_/A sky130_fd_sc_hd__inv_2
XANTENNA__15070__D _15069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _17260_/A _17247_/X VGND VGND VPWR VPWR _17336_/X sky130_fd_sc_hd__or2_4
XANTENNA__19120__A _19106_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14548_ _14548_/A VGND VGND VPWR VPWR _14548_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17267_ _17346_/B _17231_/X VGND VGND VPWR VPWR _17267_/X sky130_fd_sc_hd__and2_4
X_14479_ _14478_/Y _14476_/X _14414_/X _14476_/X VGND VGND VPWR VPWR _14479_/X sky130_fd_sc_hd__a2bb2o_4
X_19006_ _19004_/Y _19005_/X _18961_/X _19005_/X VGND VGND VPWR VPWR _23879_/D sky130_fd_sc_hd__a2bb2o_4
X_16218_ _16216_/Y _16212_/X _15959_/X _16217_/X VGND VGND VPWR VPWR _16218_/X sky130_fd_sc_hd__a2bb2o_4
X_17198_ _22478_/A _17196_/A _16342_/Y _17350_/A VGND VGND VPWR VPWR _17201_/C sky130_fd_sc_hd__o22a_4
XFILLER_122_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16149_ _22395_/A VGND VGND VPWR VPWR _16149_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18598__A2_N _18789_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15873__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19908_ _23564_/Q VGND VGND VPWR VPWR _19908_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19064__B1 _19018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19839_ _19838_/Y _19836_/X _19797_/X _19836_/X VGND VGND VPWR VPWR _19839_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22850_ _22792_/A VGND VGND VPWR VPWR _22850_/X sky130_fd_sc_hd__buf_2
XFILLER_83_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23163__A2 _22988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21801_ _21670_/A _21801_/B VGND VGND VPWR VPWR _21801_/X sky130_fd_sc_hd__or2_4
X_22781_ _22779_/X _22780_/X _22440_/C VGND VGND VPWR VPWR _22781_/X sky130_fd_sc_hd__or3_4
XANTENNA__17378__B1 _17271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24537__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14439__A _25123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21732_ _16785_/Y _22835_/A VGND VGND VPWR VPWR _21732_/X sky130_fd_sc_hd__and2_4
X_24520_ _24555_/CLK _16578_/X HRESETn VGND VGND VPWR VPWR _24520_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_33_0_HCLK clkbuf_7_16_0_HCLK/X VGND VGND VPWR VPWR _23832_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12239__A1_N _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16050__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_96_0_HCLK clkbuf_7_48_0_HCLK/X VGND VGND VPWR VPWR _24362_/CLK sky130_fd_sc_hd__clkbuf_1
X_21663_ _21663_/A VGND VGND VPWR VPWR _21664_/A sky130_fd_sc_hd__buf_2
X_24451_ _25016_/CLK _24451_/D HRESETn VGND VGND VPWR VPWR _24451_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20614_ _17389_/A _17388_/X VGND VGND VPWR VPWR _20615_/B sky130_fd_sc_hd__nand2_4
X_23402_ _23580_/CLK _23402_/D VGND VGND VPWR VPWR _23402_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22674__A1 _21095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24382_ _24391_/CLK _17089_/Y HRESETn VGND VGND VPWR VPWR _24382_/Q sky130_fd_sc_hd__dfrtp_4
X_21594_ _21245_/A VGND VGND VPWR VPWR _21595_/A sky130_fd_sc_hd__buf_2
XFILLER_123_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22806__D _22806_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23333_ _23333_/A _23333_/B VGND VGND VPWR VPWR _24061_/D sky130_fd_sc_hd__or2_4
X_20545_ _20544_/X VGND VGND VPWR VPWR _23933_/D sky130_fd_sc_hd__inv_2
XFILLER_71_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23264_ _16092_/Y _22551_/X _22843_/X _11748_/Y _22846_/X VGND VGND VPWR VPWR _23264_/X
+ sky130_fd_sc_hd__o32a_4
X_20476_ _20476_/A VGND VGND VPWR VPWR _20486_/B sky130_fd_sc_hd__inv_2
XFILLER_10_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25396__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22215_ _21595_/A _22215_/B VGND VGND VPWR VPWR _22215_/X sky130_fd_sc_hd__or2_4
X_25003_ _25001_/CLK _25003_/D HRESETn VGND VGND VPWR VPWR _14915_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25325__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23195_ _15570_/Y _22872_/B VGND VGND VPWR VPWR _23195_/X sky130_fd_sc_hd__and2_4
XFILLER_105_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22146_ _22146_/A _22145_/X VGND VGND VPWR VPWR _22146_/X sky130_fd_sc_hd__and2_4
XANTENNA__12807__A1_N _22660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22077_ _22055_/X _20174_/Y VGND VGND VPWR VPWR _22077_/X sky130_fd_sc_hd__or2_4
XFILLER_86_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15734__A1_N _12584_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21028_ _21028_/A VGND VGND VPWR VPWR _21112_/B sky130_fd_sc_hd__buf_2
XFILLER_0_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23139__C1 _23138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16829__A _24415_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18661__A1_N _16616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13850_ _23990_/Q VGND VGND VPWR VPWR _13850_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24960__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12801_ _22706_/A VGND VGND VPWR VPWR _12849_/B sky130_fd_sc_hd__inv_2
XFILLER_90_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13781_ _13780_/X VGND VGND VPWR VPWR _13782_/A sky130_fd_sc_hd__inv_2
XFILLER_16_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24278__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22979_ _23114_/A _22979_/B _22979_/C _22978_/X VGND VGND VPWR VPWR _22979_/X sky130_fd_sc_hd__or4_4
XFILLER_43_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15520_ _15519_/Y _15517_/X HADDR[11] _15517_/X VGND VGND VPWR VPWR _15520_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12732_ _12730_/Y _12731_/X _12721_/X VGND VGND VPWR VPWR _25391_/D sky130_fd_sc_hd__and3_4
XFILLER_71_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24718_ _24345_/CLK _16038_/X HRESETn VGND VGND VPWR VPWR _16037_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16041__B1 _11804_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21470__A _17706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15451_ _13901_/X _15449_/X _15446_/X _13899_/X _15444_/X VGND VGND VPWR VPWR _15451_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_31_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12663_ _12662_/X VGND VGND VPWR VPWR _25410_/D sky130_fd_sc_hd__inv_2
XFILLER_93_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24649_ _24649_/CLK _16229_/X HRESETn VGND VGND VPWR VPWR _22733_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_31_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _20596_/A VGND VGND VPWR VPWR _20592_/A sky130_fd_sc_hd__inv_2
XFILLER_106_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _18202_/A _18166_/X _18170_/C VGND VGND VPWR VPWR _18178_/B sky130_fd_sc_hd__or3_4
Xclkbuf_5_4_0_HCLK clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ _15382_/A _15382_/B VGND VGND VPWR VPWR _15384_/B sky130_fd_sc_hd__or2_4
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _12606_/A _12582_/Y _12616_/B _24846_/Q VGND VGND VPWR VPWR _12598_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20086__A _20095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ _17120_/X VGND VGND VPWR VPWR _17121_/Y sky130_fd_sc_hd__inv_2
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14333_ _12163_/A _12157_/X VGND VGND VPWR VPWR _14333_/X sky130_fd_sc_hd__or2_4
XFILLER_7_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052_ _24391_/Q _17053_/B VGND VGND VPWR VPWR _17052_/X sky130_fd_sc_hd__or2_4
X_14264_ _14271_/A VGND VGND VPWR VPWR _14264_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16003_ _16002_/X VGND VGND VPWR VPWR _16003_/X sky130_fd_sc_hd__buf_2
X_13215_ _13457_/A _13211_/X _13215_/C VGND VGND VPWR VPWR _13215_/X sky130_fd_sc_hd__and3_4
XFILLER_100_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25066__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14195_ _14195_/A _14195_/B VGND VGND VPWR VPWR _14210_/B sky130_fd_sc_hd__or2_4
XFILLER_100_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13146_ _24190_/Q VGND VGND VPWR VPWR _13234_/A sky130_fd_sc_hd__buf_2
XFILLER_98_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13077_ _12347_/Y _13071_/X _13073_/Y _13031_/X VGND VGND VPWR VPWR _13077_/X sky130_fd_sc_hd__a211o_4
X_17954_ _14648_/X _17952_/X _17954_/C VGND VGND VPWR VPWR _17954_/X sky130_fd_sc_hd__and3_4
XFILLER_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19046__B1 _18997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12028_ _12028_/A VGND VGND VPWR VPWR _12034_/A sky130_fd_sc_hd__inv_2
X_16905_ _24263_/Q VGND VGND VPWR VPWR _17758_/A sky130_fd_sc_hd__inv_2
XANTENNA__17057__C1 _17056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17885_ _21048_/A _17885_/B VGND VGND VPWR VPWR _17885_/X sky130_fd_sc_hd__or2_4
XFILLER_39_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16836_ _24412_/Q VGND VGND VPWR VPWR _16836_/Y sky130_fd_sc_hd__inv_2
X_19624_ _19624_/A VGND VGND VPWR VPWR _21811_/B sky130_fd_sc_hd__inv_2
XFILLER_19_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19555_ _19555_/A VGND VGND VPWR VPWR _19555_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16767_ _24445_/Q VGND VGND VPWR VPWR _16767_/Y sky130_fd_sc_hd__inv_2
X_13979_ _25219_/Q VGND VGND VPWR VPWR _13980_/A sky130_fd_sc_hd__buf_2
XFILLER_93_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24630__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18506_ _18821_/B _18506_/B _18505_/X VGND VGND VPWR VPWR _18507_/A sky130_fd_sc_hd__or3_4
X_15718_ _15721_/A VGND VGND VPWR VPWR _15718_/X sky130_fd_sc_hd__buf_2
X_19486_ _21483_/B _19483_/X _11955_/X _19483_/X VGND VGND VPWR VPWR _23710_/D sky130_fd_sc_hd__a2bb2o_4
X_16698_ _16697_/Y _16695_/X _16600_/X _16695_/X VGND VGND VPWR VPWR _24475_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16032__B1 _15964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22476__A _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18437_ _16209_/Y _24167_/Q _22539_/A _18566_/A VGND VGND VPWR VPWR _18444_/A sky130_fd_sc_hd__a2bb2o_4
X_15649_ _15649_/A VGND VGND VPWR VPWR _15843_/A sky130_fd_sc_hd__buf_2
XANTENNA__22105__B1 _21306_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18368_ _18367_/Y _18355_/Y _18365_/A _18355_/A VGND VGND VPWR VPWR _18368_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22656__A1 _15709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22656__B2 _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17319_ _17254_/C _17323_/B _17318_/Y VGND VGND VPWR VPWR _17319_/X sky130_fd_sc_hd__o21a_4
X_18299_ _18298_/X VGND VGND VPWR VPWR _18299_/X sky130_fd_sc_hd__buf_2
X_20330_ _20317_/X _19586_/D _18254_/X _21977_/B _20326_/A VGND VGND VPWR VPWR _23407_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_122_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23100__A _23100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20261_ _23433_/Q VGND VGND VPWR VPWR _21903_/B sky130_fd_sc_hd__inv_2
X_22000_ _11677_/A _22727_/B _21504_/B _21999_/Y VGND VGND VPWR VPWR _22000_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16099__B1 _15944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21092__B1 _22664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17835__A1 _17755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20192_ _22357_/B _20191_/X _19777_/A _20191_/X VGND VGND VPWR VPWR _23460_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13537__A1_N _13536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24789__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23951_ _25137_/CLK _23951_/D HRESETn VGND VGND VPWR VPWR _23951_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24718__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15553__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22902_ _22902_/A _22864_/X VGND VGND VPWR VPWR _22902_/X sky130_fd_sc_hd__or2_4
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23882_ _23884_/CLK _23882_/D VGND VGND VPWR VPWR _18995_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_99_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_4_0_HCLK_A clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22833_ _21066_/A VGND VGND VPWR VPWR _22833_/X sky130_fd_sc_hd__buf_2
XANTENNA__21147__A1 _21350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24371__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12178__A1_N _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12832__B1 _12819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24300__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22764_ _22764_/A VGND VGND VPWR VPWR _22897_/A sky130_fd_sc_hd__buf_2
XANTENNA__16023__B1 _15955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24503_ _24502_/CLK _24503_/D HRESETn VGND VGND VPWR VPWR _16620_/A sky130_fd_sc_hd__dfrtp_4
X_21715_ _17429_/Y _21549_/B VGND VGND VPWR VPWR _21715_/Y sky130_fd_sc_hd__nor2_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25483_ _23689_/CLK _11988_/X HRESETn VGND VGND VPWR VPWR _11654_/B sky130_fd_sc_hd__dfrtp_4
X_22695_ _24447_/Q _22695_/B _22695_/C VGND VGND VPWR VPWR _22695_/X sky130_fd_sc_hd__and3_4
XFILLER_129_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16384__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21646_ _21634_/Y _21645_/Y _13784_/C VGND VGND VPWR VPWR _21646_/X sky130_fd_sc_hd__o21a_4
X_24434_ _24596_/CLK _24434_/D HRESETn VGND VGND VPWR VPWR _24434_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20658__B1 _17401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21577_ _22441_/A _21572_/X _22444_/A _21576_/X VGND VGND VPWR VPWR _21578_/B sky130_fd_sc_hd__o22a_4
XANTENNA__25506__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24365_ _24368_/CLK _24365_/D HRESETn VGND VGND VPWR VPWR _16994_/A sky130_fd_sc_hd__dfrtp_4
X_20528_ _20427_/C _20433_/X _20497_/X VGND VGND VPWR VPWR _24077_/D sky130_fd_sc_hd__a21o_4
X_23316_ _25451_/Q _21064_/X _23314_/X _23315_/X _22440_/C VGND VGND VPWR VPWR _23316_/X
+ sky130_fd_sc_hd__a2111o_4
X_24296_ _25433_/CLK _17642_/X HRESETn VGND VGND VPWR VPWR _24296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20459_ _25140_/Q _20459_/B _20457_/D VGND VGND VPWR VPWR _20459_/X sky130_fd_sc_hd__and3_4
XFILLER_84_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23247_ _23247_/A _22810_/X _22812_/C VGND VGND VPWR VPWR _23247_/X sky130_fd_sc_hd__and3_4
X_13000_ _12306_/Y _12999_/X VGND VGND VPWR VPWR _13001_/D sky130_fd_sc_hd__or2_4
XANTENNA__11975__B _11970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23178_ _23178_/A _23269_/B VGND VGND VPWR VPWR _23178_/X sky130_fd_sc_hd__or2_4
XFILLER_122_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15837__B1 _24811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22129_ _21416_/A VGND VGND VPWR VPWR _22130_/C sky130_fd_sc_hd__buf_2
XANTENNA__13248__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19028__B1 _18977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21465__A _21465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14951_ _14943_/X _14946_/X _14951_/C _14950_/X VGND VGND VPWR VPWR _14951_/X sky130_fd_sc_hd__or4_4
XANTENNA__24459__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13902_ _13901_/X VGND VGND VPWR VPWR _13905_/B sky130_fd_sc_hd__inv_2
X_17670_ _17574_/Y _17673_/B _17590_/X VGND VGND VPWR VPWR _17670_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14882_ _14872_/B _14880_/Y _14828_/X _14881_/Y _14831_/A VGND VGND VPWR VPWR _14882_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16262__B1 _15474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23127__A2 _22988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16621_ _16620_/Y _16545_/A _16266_/X _16545_/A VGND VGND VPWR VPWR _24503_/D sky130_fd_sc_hd__a2bb2o_4
X_13833_ _13821_/A VGND VGND VPWR VPWR _13833_/X sky130_fd_sc_hd__buf_2
XANTENNA__21138__A1 _13789_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19340_ _19338_/Y _19334_/X _19294_/X _19339_/X VGND VGND VPWR VPWR _23762_/D sky130_fd_sc_hd__a2bb2o_4
X_16552_ _16549_/Y _16545_/X _16380_/X _16551_/X VGND VGND VPWR VPWR _16552_/X sky130_fd_sc_hd__a2bb2o_4
X_13764_ _13746_/A _13760_/X _13762_/X _14703_/A VGND VGND VPWR VPWR _13764_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12823__B1 _25375_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24041__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15503_ _15503_/A VGND VGND VPWR VPWR _15503_/Y sky130_fd_sc_hd__inv_2
X_12715_ _12698_/A _12712_/B _12714_/Y VGND VGND VPWR VPWR _25397_/D sky130_fd_sc_hd__and3_4
X_19271_ _19278_/A VGND VGND VPWR VPWR _19271_/X sky130_fd_sc_hd__buf_2
X_16483_ _24556_/Q VGND VGND VPWR VPWR _16483_/Y sky130_fd_sc_hd__inv_2
X_13695_ _13695_/A _13695_/B VGND VGND VPWR VPWR _13695_/X sky130_fd_sc_hd__and2_4
XANTENNA__14807__A _14807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18222_ _18046_/A _18222_/B VGND VGND VPWR VPWR _18222_/X sky130_fd_sc_hd__or2_4
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15434_ _15452_/A VGND VGND VPWR VPWR _15434_/X sky130_fd_sc_hd__buf_2
XFILLER_62_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16725__C _22574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12646_ _12657_/A _12644_/X _12645_/X VGND VGND VPWR VPWR _12646_/X sky130_fd_sc_hd__and3_4
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18153_ _18185_/A _18153_/B _18153_/C VGND VGND VPWR VPWR _18161_/B sky130_fd_sc_hd__or3_4
XANTENNA__19503__B2 _19500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15365_ _15365_/A _15365_/B VGND VGND VPWR VPWR _15369_/B sky130_fd_sc_hd__or2_4
XANTENNA__25247__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12577_ _12576_/Y _24857_/Q _12576_/Y _24857_/Q VGND VGND VPWR VPWR _12578_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17104_ _16972_/Y _17108_/B _17103_/Y VGND VGND VPWR VPWR _17104_/X sky130_fd_sc_hd__o21a_4
X_14316_ _14306_/X _14315_/X _13484_/A _14311_/X VGND VGND VPWR VPWR _25162_/D sky130_fd_sc_hd__o22a_4
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18084_ _18046_/A _19000_/A VGND VGND VPWR VPWR _18085_/C sky130_fd_sc_hd__or2_4
X_15296_ _15296_/A _15365_/A _15139_/Y _15130_/Y VGND VGND VPWR VPWR _15296_/X sky130_fd_sc_hd__or4_4
XANTENNA__17837__B _17751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17035_ _17035_/A _17007_/Y _17034_/X VGND VGND VPWR VPWR _17047_/A sky130_fd_sc_hd__or3_4
X_14247_ _13886_/X _15441_/A _20490_/A VGND VGND VPWR VPWR _14247_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__18014__A _18010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14178_ _14173_/A _14173_/B _14173_/Y VGND VGND VPWR VPWR _14178_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__15828__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13129_ _13129_/A _13129_/B _20717_/A _20712_/A VGND VGND VPWR VPWR _13130_/B sky130_fd_sc_hd__or4_4
XANTENNA__19019__B1 _19018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18986_ _23884_/Q VGND VGND VPWR VPWR _18986_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24882__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17937_ _17955_/A _19126_/A VGND VGND VPWR VPWR _17939_/B sky130_fd_sc_hd__or2_4
XANTENNA__24811__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17868_ _16911_/Y _17867_/X _16955_/X VGND VGND VPWR VPWR _17868_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_61_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17291__C _17346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24129__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19607_ _19606_/Y _19602_/X _19420_/X _19587_/X VGND VGND VPWR VPWR _23669_/D sky130_fd_sc_hd__a2bb2o_4
X_16819_ _16807_/A VGND VGND VPWR VPWR _16819_/X sky130_fd_sc_hd__buf_2
X_17799_ _16909_/Y _17794_/B _17780_/X _17795_/Y VGND VGND VPWR VPWR _17799_/X sky130_fd_sc_hd__a211o_4
XFILLER_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19538_ _19538_/A VGND VGND VPWR VPWR _19538_/X sky130_fd_sc_hd__buf_2
XANTENNA__12814__B1 _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12530__A2_N _24842_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19469_ _18275_/X _20338_/B _19888_/C VGND VGND VPWR VPWR _19469_/X sky130_fd_sc_hd__or3_4
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21500_ _21495_/X _21499_/X _11683_/Y _21495_/X VGND VGND VPWR VPWR _21500_/X sky130_fd_sc_hd__a2bb2o_4
X_22480_ _21111_/X VGND VGND VPWR VPWR _22480_/X sky130_fd_sc_hd__buf_2
XANTENNA__14436__B _18895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21431_ _22963_/A VGND VGND VPWR VPWR _23271_/A sky130_fd_sc_hd__buf_2
XFILLER_124_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_107_0_HCLK clkbuf_7_53_0_HCLK/X VGND VGND VPWR VPWR _24600_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24150_ _24159_/CLK _24150_/D HRESETn VGND VGND VPWR VPWR _18581_/A sky130_fd_sc_hd__dfrtp_4
X_21362_ _19582_/X VGND VGND VPWR VPWR _21362_/X sky130_fd_sc_hd__buf_2
XFILLER_135_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20313_ _23413_/Q VGND VGND VPWR VPWR _20313_/Y sky130_fd_sc_hd__inv_2
X_23101_ _24797_/Q _23101_/B VGND VGND VPWR VPWR _23101_/X sky130_fd_sc_hd__or2_4
X_24081_ _23995_/CLK _20460_/X HRESETn VGND VGND VPWR VPWR _20444_/A sky130_fd_sc_hd__dfrtp_4
X_21293_ _21293_/A VGND VGND VPWR VPWR _21293_/X sky130_fd_sc_hd__buf_2
XANTENNA__14452__A _14381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23032_ _22759_/X _23031_/X _22854_/X _24830_/Q _22761_/X VGND VGND VPWR VPWR _23033_/B
+ sky130_fd_sc_hd__a32o_4
X_20244_ _13373_/B VGND VGND VPWR VPWR _20244_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20175_ _20182_/A VGND VGND VPWR VPWR _20175_/X sky130_fd_sc_hd__buf_2
XFILLER_88_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16492__B1 _16405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24552__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24983_ _24984_/CLK _15359_/Y HRESETn VGND VGND VPWR VPWR _24983_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23934_ _25122_/CLK _20551_/Y HRESETn VGND VGND VPWR VPWR _23934_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23865_ _25485_/CLK _23865_/D VGND VGND VPWR VPWR _19047_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_84_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22816_ _22816_/A _22394_/X _22493_/B VGND VGND VPWR VPWR _22816_/X sky130_fd_sc_hd__and3_4
XANTENNA__21732__B _22835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23796_ _24398_/CLK _23796_/D VGND VGND VPWR VPWR _23796_/Q sky130_fd_sc_hd__dfxtp_4
X_25535_ _24267_/CLK _25535_/D HRESETn VGND VGND VPWR VPWR _11753_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_77_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22747_ _15599_/Y _22747_/B VGND VGND VPWR VPWR _22747_/X sky130_fd_sc_hd__and2_4
XFILLER_25_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12500_ _12264_/X _12499_/X _12394_/X VGND VGND VPWR VPWR _12500_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_38_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13480_ _13479_/Y _13477_/X _11838_/X _13477_/X VGND VGND VPWR VPWR _13480_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_66_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_66_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_25466_ _24097_/CLK _12091_/X HRESETn VGND VGND VPWR VPWR _12090_/A sky130_fd_sc_hd__dfrtp_4
X_22678_ _21106_/X _22676_/X _21211_/X _22677_/X VGND VGND VPWR VPWR _22679_/B sky130_fd_sc_hd__o22a_4
X_12431_ _12249_/X _12238_/X _12430_/X VGND VGND VPWR VPWR _12432_/B sky130_fd_sc_hd__or3_4
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24417_ _24462_/CLK _16826_/X HRESETn VGND VGND VPWR VPWR _16823_/A sky130_fd_sc_hd__dfrtp_4
X_21629_ _21629_/A _21629_/B VGND VGND VPWR VPWR _21631_/B sky130_fd_sc_hd__or2_4
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25340__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25397_ _25397_/CLK _25397_/D HRESETn VGND VGND VPWR VPWR _25397_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15150_ _24983_/Q VGND VGND VPWR VPWR _15298_/B sky130_fd_sc_hd__inv_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12362_ _12999_/B _12368_/A _12992_/A _12305_/Y VGND VGND VPWR VPWR _12371_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23966__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24348_ _24330_/CLK _24348_/D HRESETn VGND VGND VPWR VPWR _22939_/A sky130_fd_sc_hd__dfrtp_4
X_14101_ _25205_/Q _14101_/B _14116_/A VGND VGND VPWR VPWR _14102_/B sky130_fd_sc_hd__or3_4
XANTENNA__11792__B1 _11791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12293_ _12292_/Y _24818_/Q _12292_/Y _24818_/Q VGND VGND VPWR VPWR _12293_/X sky130_fd_sc_hd__a2bb2o_4
X_15081_ _15080_/Y _24592_/Q _15080_/Y _24592_/Q VGND VGND VPWR VPWR _15082_/D sky130_fd_sc_hd__a2bb2o_4
X_24279_ _24278_/CLK _24279_/D HRESETn VGND VGND VPWR VPWR _17527_/A sky130_fd_sc_hd__dfrtp_4
X_14032_ _14023_/A VGND VGND VPWR VPWR _14032_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18840_ _24561_/Q _18696_/A _16537_/Y _24114_/Q VGND VGND VPWR VPWR _18843_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16078__A3 _15927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18771_ _18771_/A VGND VGND VPWR VPWR _18771_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15825__A3 _11818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15983_ _12232_/Y _15982_/X _15627_/X _15982_/X VGND VGND VPWR VPWR _24740_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16289__A _16288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24293__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17722_ _17722_/A VGND VGND VPWR VPWR _17722_/X sky130_fd_sc_hd__buf_2
X_14934_ _14934_/A VGND VGND VPWR VPWR _14934_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19421__B1 _19420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24222__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17653_ _17611_/A _17653_/B VGND VGND VPWR VPWR _17653_/X sky130_fd_sc_hd__or2_4
XANTENNA__21923__A _21944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14865_ _14880_/B _14798_/X _25031_/Q _14864_/X VGND VGND VPWR VPWR _14865_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16604_ HWDATA[8] VGND VGND VPWR VPWR _16604_/X sky130_fd_sc_hd__buf_2
XFILLER_63_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13816_ _13815_/X VGND VGND VPWR VPWR _13817_/A sky130_fd_sc_hd__inv_2
XFILLER_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17584_ _17611_/A _17597_/A _17584_/C _17583_/X VGND VGND VPWR VPWR _17585_/B sky130_fd_sc_hd__or4_4
XANTENNA__25499__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14796_ scl_oen_o_S5 _20996_/B _14796_/C VGND VGND VPWR VPWR _14807_/B sky130_fd_sc_hd__and3_4
XFILLER_17_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19323_ _19322_/Y _19318_/X _19232_/X _19318_/X VGND VGND VPWR VPWR _19323_/X sky130_fd_sc_hd__a2bb2o_4
X_16535_ _16535_/A VGND VGND VPWR VPWR _16535_/Y sky130_fd_sc_hd__inv_2
X_13747_ _13757_/A VGND VGND VPWR VPWR _13748_/C sky130_fd_sc_hd__buf_2
XANTENNA__25428__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16538__B2 _16461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18009__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19254_ _19253_/Y _19249_/X _16881_/X _19249_/X VGND VGND VPWR VPWR _23792_/D sky130_fd_sc_hd__a2bb2o_4
X_16466_ _16466_/A VGND VGND VPWR VPWR _16474_/A sky130_fd_sc_hd__buf_2
X_13678_ _13713_/A _13678_/B VGND VGND VPWR VPWR _13694_/B sky130_fd_sc_hd__or2_4
XFILLER_108_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18205_ _14646_/X _18203_/X _18205_/C VGND VGND VPWR VPWR _18205_/X sky130_fd_sc_hd__and3_4
X_15417_ _15159_/X _15415_/X VGND VGND VPWR VPWR _15417_/X sky130_fd_sc_hd__or2_4
X_12629_ _12693_/A _12602_/A VGND VGND VPWR VPWR _12629_/X sky130_fd_sc_hd__and2_4
X_19185_ _23816_/Q VGND VGND VPWR VPWR _19185_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25081__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16397_ _16396_/Y _16394_/X _16306_/X _16394_/X VGND VGND VPWR VPWR _16397_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18136_ _18104_/A _20223_/A VGND VGND VPWR VPWR _18136_/X sky130_fd_sc_hd__or2_4
XFILLER_8_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15348_ _15315_/A _15345_/B _15347_/X VGND VGND VPWR VPWR _15349_/A sky130_fd_sc_hd__or3_4
XANTENNA__25010__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18067_ _18104_/A _23449_/Q VGND VGND VPWR VPWR _18068_/C sky130_fd_sc_hd__or2_4
X_15279_ _14981_/X _15282_/B _15174_/X VGND VGND VPWR VPWR _15279_/Y sky130_fd_sc_hd__a21oi_4
X_17018_ _16990_/X _17017_/X VGND VGND VPWR VPWR _17346_/B sky130_fd_sc_hd__or2_4
XFILLER_99_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18969_ _23891_/Q VGND VGND VPWR VPWR _18969_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13616__A _17995_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21980_ _18270_/X _21967_/X _21971_/Y _21504_/B _21979_/X VGND VGND VPWR VPWR _21980_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18430__A1_N _16230_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16226__B1 _11796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22929__A _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20931_ _20931_/A _20931_/B VGND VGND VPWR VPWR _20931_/X sky130_fd_sc_hd__or2_4
XFILLER_94_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20862_ _24039_/Q _13659_/X _20861_/Y VGND VGND VPWR VPWR _20862_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23650_ _23649_/CLK _19670_/X VGND VGND VPWR VPWR _19668_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23945__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22601_ _22146_/A _22596_/X _21826_/X _22600_/Y VGND VGND VPWR VPWR _22602_/A sky130_fd_sc_hd__a211o_4
XANTENNA__18445__A1_N _16261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20793_ _20790_/Y _20791_/Y _20792_/X VGND VGND VPWR VPWR _20793_/X sky130_fd_sc_hd__o21a_4
XFILLER_22_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23581_ _23581_/CLK _19864_/X VGND VGND VPWR VPWR _23581_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17726__B1 _17722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25320_ _23377_/CLK _25320_/D HRESETn VGND VGND VPWR VPWR _25320_/Q sky130_fd_sc_hd__dfrtp_4
X_22532_ _22532_/A _22727_/B VGND VGND VPWR VPWR _22532_/X sky130_fd_sc_hd__and2_4
XFILLER_50_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25251_ _25263_/CLK _25251_/D HRESETn VGND VGND VPWR VPWR _13831_/A sky130_fd_sc_hd__dfrtp_4
X_22463_ _22434_/X _22440_/X _22447_/Y _22462_/X VGND VGND VPWR VPWR HRDATA[8] sky130_fd_sc_hd__a211o_4
XFILLER_72_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22383__B _22301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24202_ _24290_/CLK _18297_/X HRESETn VGND VGND VPWR VPWR _24202_/Q sky130_fd_sc_hd__dfrtp_4
X_21414_ _21414_/A _21073_/B VGND VGND VPWR VPWR _21414_/X sky130_fd_sc_hd__or2_4
X_22394_ _22836_/B VGND VGND VPWR VPWR _22394_/X sky130_fd_sc_hd__buf_2
X_25182_ _24148_/CLK _14240_/X HRESETn VGND VGND VPWR VPWR _14238_/A sky130_fd_sc_hd__dfstp_4
X_21345_ _13514_/Y _12096_/X _12043_/Y _16453_/B VGND VGND VPWR VPWR _21345_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24133_ _24133_/CLK _18752_/Y HRESETn VGND VGND VPWR VPWR _24133_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21276_ _15551_/B VGND VGND VPWR VPWR _22827_/A sky130_fd_sc_hd__buf_2
X_24064_ _24957_/CLK _24064_/D HRESETn VGND VGND VPWR VPWR HREADYOUT sky130_fd_sc_hd__dfstp_4
XANTENNA__23498__CLK _23498_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24733__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_HCLK clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_20227_ _20226_/Y _20224_/X _18267_/X _20224_/X VGND VGND VPWR VPWR _23446_/D sky130_fd_sc_hd__a2bb2o_4
X_23015_ _16666_/Y _22824_/X _15583_/Y _22827_/X VGND VGND VPWR VPWR _23015_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19651__B1 _19599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20158_ _23472_/Q VGND VGND VPWR VPWR _20158_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15807__A3 _15729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12980_ _12980_/A VGND VGND VPWR VPWR _12980_/Y sky130_fd_sc_hd__inv_2
X_20089_ _20089_/A VGND VGND VPWR VPWR _20089_/X sky130_fd_sc_hd__buf_2
XANTENNA__12430__A _12430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24966_ _24977_/CLK _24966_/D HRESETn VGND VGND VPWR VPWR _24966_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_94_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11931_ _11929_/Y _11926_/X _11930_/X _11926_/X VGND VGND VPWR VPWR _11931_/X sky130_fd_sc_hd__a2bb2o_4
X_23917_ _23959_/CLK _20529_/X HRESETn VGND VGND VPWR VPWR _23917_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24897_ _24868_/CLK _15596_/X HRESETn VGND VGND VPWR VPWR _15595_/A sky130_fd_sc_hd__dfrtp_4
X_14650_ _17975_/A VGND VGND VPWR VPWR _18010_/A sky130_fd_sc_hd__buf_2
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11862_ _11862_/A VGND VGND VPWR VPWR _11862_/X sky130_fd_sc_hd__buf_2
XFILLER_72_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23848_ _23847_/CLK _23848_/D VGND VGND VPWR VPWR _19095_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_45_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13601_ _19038_/D VGND VGND VPWR VPWR _13633_/B sky130_fd_sc_hd__buf_2
X_14581_ _13570_/Y _14581_/B VGND VGND VPWR VPWR _14581_/X sky130_fd_sc_hd__or2_4
XANTENNA__25521__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11793_ _25523_/Q VGND VGND VPWR VPWR _11793_/Y sky130_fd_sc_hd__inv_2
X_23779_ _23618_/CLK _23779_/D VGND VGND VPWR VPWR _13240_/B sky130_fd_sc_hd__dfxtp_4
X_16320_ _22816_/A VGND VGND VPWR VPWR _16320_/Y sky130_fd_sc_hd__inv_2
X_13532_ _13532_/A VGND VGND VPWR VPWR SSn_S2 sky130_fd_sc_hd__inv_2
X_25518_ _25514_/CLK _25518_/D HRESETn VGND VGND VPWR VPWR _25518_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22574__A _22574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17193__B2 _17254_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16251_ _22294_/A VGND VGND VPWR VPWR _16251_/Y sky130_fd_sc_hd__inv_2
X_13463_ _13199_/Y _13447_/X _13462_/X _25314_/Q _11964_/X VGND VGND VPWR VPWR _13463_/X
+ sky130_fd_sc_hd__o32a_4
X_25449_ _25449_/CLK _12401_/X HRESETn VGND VGND VPWR VPWR _12399_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16572__A _24522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22293__B _22293_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15202_ _15193_/B VGND VGND VPWR VPWR _15203_/B sky130_fd_sc_hd__inv_2
X_12414_ _12252_/Y _12288_/X _12382_/X VGND VGND VPWR VPWR _12414_/X sky130_fd_sc_hd__or3_4
X_16182_ _16449_/A VGND VGND VPWR VPWR _22444_/A sky130_fd_sc_hd__buf_2
X_13394_ _13426_/A _23615_/Q VGND VGND VPWR VPWR _13396_/B sky130_fd_sc_hd__or2_4
XFILLER_16_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11765__B1 _11764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_153_0_HCLK clkbuf_7_76_0_HCLK/X VGND VGND VPWR VPWR _25514_/CLK sky130_fd_sc_hd__clkbuf_1
X_15133_ _15382_/A VGND VGND VPWR VPWR _15133_/Y sky130_fd_sc_hd__inv_2
X_12345_ _12345_/A VGND VGND VPWR VPWR _12345_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12605__A _12665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15064_ _15064_/A _15267_/A _15064_/C _15063_/X VGND VGND VPWR VPWR _15209_/C sky130_fd_sc_hd__or4_4
X_19941_ _21796_/B _19936_/X _19625_/X _19936_/X VGND VGND VPWR VPWR _19941_/X sky130_fd_sc_hd__a2bb2o_4
X_12276_ _25448_/Q VGND VGND VPWR VPWR _12385_/B sky130_fd_sc_hd__inv_2
XANTENNA__24474__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14015_ _13984_/X _13995_/X _14006_/X _14538_/D VGND VGND VPWR VPWR _14015_/X sky130_fd_sc_hd__a211o_4
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19872_ _23578_/Q VGND VGND VPWR VPWR _19872_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24403__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16456__B1 _16366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18823_ pwm_S7 VGND VGND VPWR VPWR _18823_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16233__A1_N _16230_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15966_ _15795_/A VGND VGND VPWR VPWR _15966_/X sky130_fd_sc_hd__buf_2
X_18754_ _18626_/Y _18759_/B _18707_/X VGND VGND VPWR VPWR _18754_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16208__B1 _11771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21201__B1 _23342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14917_ _14915_/A _24409_/Q _15063_/B _14916_/Y VGND VGND VPWR VPWR _14917_/X sky130_fd_sc_hd__o22a_4
X_17705_ _21194_/A VGND VGND VPWR VPWR _17706_/A sky130_fd_sc_hd__buf_2
XFILLER_82_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15897_ _11821_/X VGND VGND VPWR VPWR _15897_/X sky130_fd_sc_hd__buf_2
X_18685_ _24126_/Q VGND VGND VPWR VPWR _18692_/A sky130_fd_sc_hd__inv_2
XFILLER_64_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14848_ _14845_/X _14847_/Y _14238_/A _14845_/X VGND VGND VPWR VPWR _14848_/X sky130_fd_sc_hd__a2bb2o_4
X_17636_ _17521_/Y _17525_/Y _17564_/Y _17645_/B VGND VGND VPWR VPWR _17642_/B sky130_fd_sc_hd__or4_4
XFILLER_24_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16248__A1_N _16246_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22187__C _22179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17567_ _17567_/A _17564_/Y _17565_/Y _17567_/D VGND VGND VPWR VPWR _17567_/X sky130_fd_sc_hd__or4_4
XANTENNA__25262__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14779_ _25046_/Q _14783_/A _14772_/X _14778_/Y VGND VGND VPWR VPWR _25046_/D sky130_fd_sc_hd__o22a_4
XFILLER_90_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12245__B2 _24758_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16518_ _16518_/A VGND VGND VPWR VPWR _16518_/Y sky130_fd_sc_hd__inv_2
X_19306_ _13451_/B VGND VGND VPWR VPWR _19306_/Y sky130_fd_sc_hd__inv_2
X_17498_ _11793_/Y _24294_/Q _11793_/Y _24294_/Q VGND VGND VPWR VPWR _17505_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16449_ _16449_/A VGND VGND VPWR VPWR _22088_/A sky130_fd_sc_hd__inv_2
X_19237_ _13404_/B VGND VGND VPWR VPWR _19237_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21268__B1 _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19168_ _19166_/Y _19167_/X _19077_/X _19167_/X VGND VGND VPWR VPWR _23823_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18119_ _18215_/A _23880_/Q VGND VGND VPWR VPWR _18120_/C sky130_fd_sc_hd__or2_4
XANTENNA__19793__A _19793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19099_ _19097_/Y _19098_/X _16885_/X _19098_/X VGND VGND VPWR VPWR _19099_/X sky130_fd_sc_hd__a2bb2o_4
X_21130_ _12054_/X _21128_/X _13468_/X _21129_/X VGND VGND VPWR VPWR _21130_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21061_ _21045_/X _21048_/X _21060_/X VGND VGND VPWR VPWR _21061_/X sky130_fd_sc_hd__and3_4
XANTENNA__24144__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18202__A _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20012_ _21793_/B _20007_/X _19988_/X _20007_/X VGND VGND VPWR VPWR _20012_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_28_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24820_ _24821_/CLK _15822_/X HRESETn VGND VGND VPWR VPWR _24820_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22659__A _22659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24751_ _24766_/CLK _15968_/X HRESETn VGND VGND VPWR VPWR _24751_/Q sky130_fd_sc_hd__dfrtp_4
X_21963_ _22385_/A _22220_/A _21963_/C _21963_/D VGND VGND VPWR VPWR _21963_/X sky130_fd_sc_hd__or4_4
XANTENNA__21743__A1 _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23702_ _23398_/CLK _19510_/X VGND VGND VPWR VPWR _23702_/Q sky130_fd_sc_hd__dfxtp_4
X_20914_ _20909_/X _20912_/X _24487_/Q _20913_/X VGND VGND VPWR VPWR _24050_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24682_ _24682_/CLK _16132_/X HRESETn VGND VGND VPWR VPWR _16130_/A sky130_fd_sc_hd__dfrtp_4
X_21894_ _21889_/X _21893_/X _14749_/A VGND VGND VPWR VPWR _21894_/X sky130_fd_sc_hd__o21a_4
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23633_ _23649_/CLK _23633_/D VGND VGND VPWR VPWR _23633_/Q sky130_fd_sc_hd__dfxtp_4
X_20845_ _20816_/X VGND VGND VPWR VPWR _20845_/X sky130_fd_sc_hd__buf_2
XANTENNA__22299__A2 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12236__B2 _24747_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23564_ _23562_/CLK _23564_/D VGND VGND VPWR VPWR _23564_/Q sky130_fd_sc_hd__dfxtp_4
X_20776_ _20772_/C _13120_/X VGND VGND VPWR VPWR _20776_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22394__A _22836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25303_ _25290_/CLK _13499_/X HRESETn VGND VGND VPWR VPWR _12023_/A sky130_fd_sc_hd__dfrtp_4
X_22515_ _21024_/A _21741_/A VGND VGND VPWR VPWR _22515_/X sky130_fd_sc_hd__or2_4
XANTENNA__23248__A1 _24732_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23495_ _23478_/CLK _20097_/X VGND VGND VPWR VPWR _20094_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24985__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25234_ _24151_/CLK _25234_/D HRESETn VGND VGND VPWR VPWR _21716_/A sky130_fd_sc_hd__dfrtp_4
X_22446_ _22441_/X _22443_/X _22444_/X _22445_/X VGND VGND VPWR VPWR _22447_/B sky130_fd_sc_hd__o22a_4
XFILLER_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11747__B1 _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24914__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25165_ _25309_/CLK _25165_/D HRESETn VGND VGND VPWR VPWR MSO_S2 sky130_fd_sc_hd__dfrtp_4
X_22377_ _22070_/X _19843_/Y _22078_/X VGND VGND VPWR VPWR _22377_/X sky130_fd_sc_hd__o21a_4
XFILLER_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_226_0_HCLK clkbuf_8_227_0_HCLK/A VGND VGND VPWR VPWR _24792_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20482__A1 _14205_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12130_ _12128_/A _12128_/B _12129_/Y VGND VGND VPWR VPWR _12130_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16686__B1 _15745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24116_ _24117_/CLK _18816_/X HRESETn VGND VGND VPWR VPWR _18681_/A sky130_fd_sc_hd__dfrtp_4
X_21328_ _16620_/A _21323_/X _15667_/A _21327_/X VGND VGND VPWR VPWR _21329_/C sky130_fd_sc_hd__a211o_4
X_25096_ _25137_/CLK _25096_/D HRESETn VGND VGND VPWR VPWR _25096_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23221__A2_N _23218_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12061_ _12060_/X VGND VGND VPWR VPWR _12061_/Y sky130_fd_sc_hd__inv_2
X_21259_ _14714_/X _21251_/X _21259_/C VGND VGND VPWR VPWR _21259_/X sky130_fd_sc_hd__or3_4
XANTENNA__22223__A2 _22727_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24047_ _24049_/CLK _24047_/D HRESETn VGND VGND VPWR VPWR _24047_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14640__A _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16438__B1 _16355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15820_ _15816_/X _15819_/X _11800_/A _24822_/Q _15817_/X VGND VGND VPWR VPWR _15820_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_38_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15751_ _15749_/X _15742_/X _15750_/X _24854_/Q _15740_/X VGND VGND VPWR VPWR _15751_/X
+ sky130_fd_sc_hd__a32o_4
X_12963_ _12833_/Y _12960_/B VGND VGND VPWR VPWR _12963_/Y sky130_fd_sc_hd__nand2_4
X_24949_ _24950_/CLK _15457_/X HRESETn VGND VGND VPWR VPWR _13895_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22931__B1 _22524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16567__A _24524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14702_ _21614_/A _14701_/X _21614_/A _14701_/X VGND VGND VPWR VPWR _14702_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15471__A _16355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11914_ _11876_/X _11916_/B VGND VGND VPWR VPWR _11914_/X sky130_fd_sc_hd__and2_4
X_18470_ _24148_/Q VGND VGND VPWR VPWR _18472_/A sky130_fd_sc_hd__inv_2
X_15682_ _15687_/A _15687_/B _15682_/C VGND VGND VPWR VPWR _15682_/X sky130_fd_sc_hd__or3_4
XFILLER_2_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12894_ _12894_/A VGND VGND VPWR VPWR _25379_/D sky130_fd_sc_hd__inv_2
X_17421_ _15623_/A VGND VGND VPWR VPWR _17421_/X sky130_fd_sc_hd__buf_2
XANTENNA__16610__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14633_ _14622_/A _14617_/Y _14632_/X _21958_/A _14622_/Y VGND VGND VPWR VPWR _25067_/D
+ sky130_fd_sc_hd__a32o_4
X_11845_ HWDATA[4] VGND VGND VPWR VPWR _15766_/A sky130_fd_sc_hd__buf_2
XFILLER_72_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17352_ _17240_/A _17352_/B VGND VGND VPWR VPWR _17354_/B sky130_fd_sc_hd__or2_4
XFILLER_54_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14564_ _13559_/Y _14601_/B VGND VGND VPWR VPWR _14564_/X sky130_fd_sc_hd__or2_4
X_11776_ _11776_/A VGND VGND VPWR VPWR _11776_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16303_ _16288_/X VGND VGND VPWR VPWR _16303_/X sky130_fd_sc_hd__buf_2
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13515_ _11862_/A VGND VGND VPWR VPWR _13515_/X sky130_fd_sc_hd__buf_2
X_17283_ _17283_/A VGND VGND VPWR VPWR _17284_/B sky130_fd_sc_hd__inv_2
X_14495_ _20428_/B VGND VGND VPWR VPWR _14495_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_36_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_73_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19022_ _23874_/Q VGND VGND VPWR VPWR _19022_/Y sky130_fd_sc_hd__inv_2
X_16234_ _24647_/Q VGND VGND VPWR VPWR _16234_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17531__A1_N _11802_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13446_ _13162_/A _13442_/X _13446_/C VGND VGND VPWR VPWR _13447_/C sky130_fd_sc_hd__or3_4
XANTENNA__24655__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16165_ _21051_/A VGND VGND VPWR VPWR _16165_/Y sky130_fd_sc_hd__inv_2
X_13377_ _13345_/A _18959_/A VGND VGND VPWR VPWR _13377_/X sky130_fd_sc_hd__or2_4
XFILLER_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15116_ _15114_/A _15115_/A _15388_/B _15115_/Y VGND VGND VPWR VPWR _15116_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16677__B1 _16408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12328_ _24836_/Q VGND VGND VPWR VPWR _12328_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16096_ _23219_/A VGND VGND VPWR VPWR _16096_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17546__A1_N _11850_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15047_ _15041_/X _15047_/B _15047_/C _15047_/D VGND VGND VPWR VPWR _15055_/C sky130_fd_sc_hd__or4_4
X_19924_ _21618_/B _19923_/X _19794_/X _19923_/X VGND VGND VPWR VPWR _19924_/X sky130_fd_sc_hd__a2bb2o_4
X_12259_ _24757_/Q VGND VGND VPWR VPWR _12259_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19855_ _21899_/B _19852_/X _19787_/X _19852_/X VGND VGND VPWR VPWR _19855_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18806_ _18782_/X _18803_/B VGND VGND VPWR VPWR _18806_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__17861__A _16918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12070__A _16453_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19786_ _19786_/A VGND VGND VPWR VPWR _21881_/B sky130_fd_sc_hd__inv_2
XFILLER_7_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16998_ _16998_/A _16998_/B _16996_/X _16997_/X VGND VGND VPWR VPWR _16998_/X sky130_fd_sc_hd__or4_4
XANTENNA__18676__B _18675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18737_ _18647_/X _18737_/B VGND VGND VPWR VPWR _18738_/C sky130_fd_sc_hd__or2_4
X_15949_ HWDATA[24] VGND VGND VPWR VPWR _15949_/X sky130_fd_sc_hd__buf_2
XANTENNA__25443__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18668_ _18668_/A _18667_/X VGND VGND VPWR VPWR _18669_/A sky130_fd_sc_hd__or2_4
XFILLER_52_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17619_ _24301_/Q _17618_/Y VGND VGND VPWR VPWR _17619_/X sky130_fd_sc_hd__or2_4
XANTENNA__12218__A1 _12399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_118_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_237_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18599_ _24144_/Q VGND VGND VPWR VPWR _18599_/X sky130_fd_sc_hd__buf_2
XFILLER_17_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20630_ _17392_/X _20630_/B _20611_/C VGND VGND VPWR VPWR _20630_/X sky130_fd_sc_hd__and3_4
XFILLER_75_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20561_ _18875_/A _18875_/B VGND VGND VPWR VPWR _20561_/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22300_ _14922_/A _21323_/X _15667_/A _22299_/X VGND VGND VPWR VPWR _22301_/C sky130_fd_sc_hd__a211o_4
XFILLER_137_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20492_ _14278_/A _20485_/B _24075_/Q VGND VGND VPWR VPWR _20494_/A sky130_fd_sc_hd__and3_4
XFILLER_30_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23280_ _23105_/X _23277_/Y _23150_/X _23279_/X VGND VGND VPWR VPWR _23280_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24396__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22942__A _22270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22231_ _22246_/A _19614_/Y VGND VGND VPWR VPWR _22231_/X sky130_fd_sc_hd__or2_4
X_22162_ _22161_/Y _21336_/A _14128_/Y _14220_/A VGND VGND VPWR VPWR _22162_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21558__A _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21113_ _21029_/X _21110_/X _21111_/X _21112_/Y VGND VGND VPWR VPWR _21114_/C sky130_fd_sc_hd__a211o_4
XFILLER_133_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15556__A _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22093_ _22701_/A _22093_/B _22093_/C VGND VGND VPWR VPWR _22093_/X sky130_fd_sc_hd__and3_4
XANTENNA__15340__B1 _15339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_56_0_HCLK clkbuf_8_57_0_HCLK/A VGND VGND VPWR VPWR _25263_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_87_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21044_ _21043_/Y VGND VGND VPWR VPWR _22146_/A sky130_fd_sc_hd__buf_2
XANTENNA__19082__B2 _19062_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23960__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24803_ _24832_/CLK _24803_/D HRESETn VGND VGND VPWR VPWR _24803_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12457__A1 _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22995_ _23133_/A _22995_/B _22995_/C VGND VGND VPWR VPWR _23002_/C sky130_fd_sc_hd__and3_4
X_24734_ _24356_/CLK _24734_/D HRESETn VGND VGND VPWR VPWR _24734_/Q sky130_fd_sc_hd__dfrtp_4
X_21946_ _21912_/X _21944_/X _21945_/X VGND VGND VPWR VPWR _21946_/X sky130_fd_sc_hd__and3_4
XANTENNA__25113__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24665_ _24654_/CLK _16188_/X HRESETn VGND VGND VPWR VPWR _23323_/A sky130_fd_sc_hd__dfrtp_4
X_21877_ _21249_/A VGND VGND VPWR VPWR _21904_/A sky130_fd_sc_hd__buf_2
XFILLER_70_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22836__B _22836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _23683_/CLK _19764_/X VGND VGND VPWR VPWR _13362_/B sky130_fd_sc_hd__dfxtp_4
X_20828_ _13655_/A VGND VGND VPWR VPWR _20828_/Y sky130_fd_sc_hd__inv_2
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24596_ _24596_/CLK _24596_/D HRESETn VGND VGND VPWR VPWR _24596_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23547_ _23388_/CLK _19955_/X VGND VGND VPWR VPWR _19954_/A sky130_fd_sc_hd__dfxtp_4
X_20759_ _20757_/Y _20754_/X _20758_/X VGND VGND VPWR VPWR _20759_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22692__A2 _22690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13260_/X _13298_/X _13299_/X VGND VGND VPWR VPWR _13300_/X sky130_fd_sc_hd__and3_4
XFILLER_13_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14280_ _15449_/A VGND VGND VPWR VPWR _14280_/X sky130_fd_sc_hd__buf_2
XANTENNA__14906__B1 _25022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23478_ _23478_/CLK _23478_/D VGND VGND VPWR VPWR _23478_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22852__A _22814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ _13143_/X _13216_/X _13231_/C VGND VGND VPWR VPWR _13231_/X sky130_fd_sc_hd__and3_4
X_25217_ _25219_/CLK _14087_/X HRESETn VGND VGND VPWR VPWR _13983_/A sky130_fd_sc_hd__dfrtp_4
X_22429_ _22429_/A VGND VGND VPWR VPWR _22714_/A sky130_fd_sc_hd__buf_2
XFILLER_40_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24066__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16850__A _16850_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16659__B1 _16300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13162_ _13162_/A VGND VGND VPWR VPWR _13162_/X sky130_fd_sc_hd__buf_2
X_25148_ _25309_/CLK _25148_/D HRESETn VGND VGND VPWR VPWR MSO_S3 sky130_fd_sc_hd__dfrtp_4
XANTENNA__15979__A1_N _12204_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12113_ _12113_/A VGND VGND VPWR VPWR _12113_/Y sky130_fd_sc_hd__inv_2
X_13093_ _13076_/A _13086_/X _13093_/C VGND VGND VPWR VPWR _25331_/D sky130_fd_sc_hd__and3_4
X_17970_ _18176_/A _17967_/X _17969_/X VGND VGND VPWR VPWR _17970_/X sky130_fd_sc_hd__and3_4
X_25079_ _25081_/CLK _14593_/X HRESETn VGND VGND VPWR VPWR _25079_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12044_ _12043_/Y _12041_/X _25475_/Q _12041_/X VGND VGND VPWR VPWR _25476_/D sky130_fd_sc_hd__a2bb2o_4
X_16921_ _21513_/A _24247_/Q _16161_/Y _16920_/Y VGND VGND VPWR VPWR _16922_/D sky130_fd_sc_hd__o22a_4
XFILLER_78_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21955__A1 _18261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21955__B2 _21636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19640_ _19636_/Y _19639_/X _19426_/X _19639_/X VGND VGND VPWR VPWR _23660_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17681__A _17624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16852_ _16442_/A VGND VGND VPWR VPWR _16852_/X sky130_fd_sc_hd__buf_2
XFILLER_93_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23157__B1 _25381_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16831__B1 _15745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15803_ _12309_/Y _15799_/X _11757_/X _15802_/X VGND VGND VPWR VPWR _24834_/D sky130_fd_sc_hd__a2bb2o_4
X_16783_ _16733_/A VGND VGND VPWR VPWR _16783_/X sky130_fd_sc_hd__buf_2
X_19571_ _23680_/Q VGND VGND VPWR VPWR _21810_/B sky130_fd_sc_hd__inv_2
XFILLER_115_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13995_ _13995_/A _13995_/B VGND VGND VPWR VPWR _13995_/X sky130_fd_sc_hd__and2_4
XFILLER_20_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21707__A1 _21275_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16297__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15734_ _12584_/Y _15732_/X _11781_/X _15732_/X VGND VGND VPWR VPWR _15734_/X sky130_fd_sc_hd__a2bb2o_4
X_18522_ _16448_/A _18478_/B VGND VGND VPWR VPWR _18523_/B sky130_fd_sc_hd__or2_4
XFILLER_98_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12946_ _25366_/Q _12945_/Y VGND VGND VPWR VPWR _12946_/X sky130_fd_sc_hd__or2_4
XFILLER_98_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15665_ _15665_/A VGND VGND VPWR VPWR _21556_/A sky130_fd_sc_hd__buf_2
X_18453_ _18772_/A VGND VGND VPWR VPWR _18521_/A sky130_fd_sc_hd__buf_2
XFILLER_60_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12877_ _12602_/A _12877_/B VGND VGND VPWR VPWR _12880_/B sky130_fd_sc_hd__or2_4
X_14616_ _14615_/Y _13638_/A _21958_/A _13637_/A VGND VGND VPWR VPWR _14616_/X sky130_fd_sc_hd__o22a_4
X_17404_ _17404_/A VGND VGND VPWR VPWR _17404_/X sky130_fd_sc_hd__buf_2
X_11828_ _11828_/A VGND VGND VPWR VPWR _11828_/Y sky130_fd_sc_hd__inv_2
X_18384_ _18377_/A VGND VGND VPWR VPWR _18384_/X sky130_fd_sc_hd__buf_2
X_15596_ _15595_/Y _15593_/X _11791_/X _15593_/X VGND VGND VPWR VPWR _15596_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24836__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17334_/X VGND VGND VPWR VPWR _24342_/D sky130_fd_sc_hd__inv_2
XANTENNA__23113__A2_N _23109_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14013_/Y _14026_/Y _14547_/C _14547_/D VGND VGND VPWR VPWR _14548_/A sky130_fd_sc_hd__or4_4
X_11759_ _25533_/Q VGND VGND VPWR VPWR _11759_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17266_ _17266_/A _17263_/X _17266_/C VGND VGND VPWR VPWR _17266_/X sky130_fd_sc_hd__and3_4
XFILLER_31_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14478_ _25107_/Q VGND VGND VPWR VPWR _14478_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16217_ _16217_/A VGND VGND VPWR VPWR _16217_/X sky130_fd_sc_hd__buf_2
X_19005_ _18988_/Y VGND VGND VPWR VPWR _19005_/X sky130_fd_sc_hd__buf_2
X_13429_ _13461_/A _13429_/B _13428_/X VGND VGND VPWR VPWR _13429_/X sky130_fd_sc_hd__or3_4
X_17197_ _17196_/Y VGND VGND VPWR VPWR _17350_/A sky130_fd_sc_hd__buf_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16148_ _16146_/Y _16144_/X _16147_/X _16144_/X VGND VGND VPWR VPWR _24676_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16079_ _16079_/A _15777_/B VGND VGND VPWR VPWR _16079_/X sky130_fd_sc_hd__or2_4
XANTENNA__19496__A2_N _19495_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14280__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19907_ _21168_/B _19902_/X _19885_/X _19902_/A VGND VGND VPWR VPWR _23565_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22738__A3 _22396_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12821__A2_N _24776_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19838_ _19838_/A VGND VGND VPWR VPWR _19838_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16822__B1 HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19769_ _19768_/Y _19766_/X _19700_/X _19766_/X VGND VGND VPWR VPWR _23614_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21800_ _21664_/A _21800_/B VGND VGND VPWR VPWR _21800_/X sky130_fd_sc_hd__or2_4
XANTENNA__17378__A1 _17244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22780_ _17253_/Y _22424_/A _12752_/A _22288_/X VGND VGND VPWR VPWR _22780_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20941__A1_N _20818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21731_ _22524_/A VGND VGND VPWR VPWR _21731_/X sky130_fd_sc_hd__buf_2
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19311__A _19310_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24450_ _25016_/CLK _24450_/D HRESETn VGND VGND VPWR VPWR _24450_/Q sky130_fd_sc_hd__dfrtp_4
X_21662_ _17728_/A VGND VGND VPWR VPWR _21681_/A sky130_fd_sc_hd__buf_2
XFILLER_127_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24577__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23401_ _23682_/CLK _20346_/X VGND VGND VPWR VPWR _20344_/A sky130_fd_sc_hd__dfxtp_4
X_20613_ _20612_/X VGND VGND VPWR VPWR _23970_/D sky130_fd_sc_hd__inv_2
XANTENNA__20134__B1 _20085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24381_ _24368_/CLK _24381_/D HRESETn VGND VGND VPWR VPWR _16967_/A sky130_fd_sc_hd__dfrtp_4
X_21593_ _21238_/X VGND VGND VPWR VPWR _21631_/A sky130_fd_sc_hd__buf_2
XFILLER_127_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22674__A2 _22672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24506__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23332_ _23313_/X _23316_/X _23320_/Y _23331_/X VGND VGND VPWR VPWR HRDATA[31] sky130_fd_sc_hd__a211o_4
X_20544_ _14444_/Y _20533_/X _14452_/X _20543_/X VGND VGND VPWR VPWR _20544_/X sky130_fd_sc_hd__a211o_4
X_23263_ _12782_/Y _22707_/X _22272_/X _12546_/Y _22844_/X VGND VGND VPWR VPWR _23263_/X
+ sky130_fd_sc_hd__o32a_4
X_20475_ _20488_/A _24075_/Q VGND VGND VPWR VPWR _20487_/A sky130_fd_sc_hd__and2_4
X_25002_ _25002_/CLK _15269_/X HRESETn VGND VGND VPWR VPWR _25002_/Q sky130_fd_sc_hd__dfrtp_4
X_22214_ _21238_/X _22212_/X _22214_/C VGND VGND VPWR VPWR _22214_/X sky130_fd_sc_hd__and3_4
XANTENNA__21634__B1 _21493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21288__A _21287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23194_ _16653_/Y _23226_/B VGND VGND VPWR VPWR _23194_/X sky130_fd_sc_hd__and2_4
XFILLER_134_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22145_ _15708_/A _22144_/X _21416_/A _25512_/Q _22929_/A VGND VGND VPWR VPWR _22145_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14190__A _16371_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22076_ _21887_/X _22076_/B VGND VGND VPWR VPWR _22076_/X sky130_fd_sc_hd__or2_4
XFILLER_82_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25365__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21027_ _21027_/A _21027_/B VGND VGND VPWR VPWR _21028_/A sky130_fd_sc_hd__or2_4
XFILLER_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12800_ _12799_/X _22623_/A _12799_/A _22623_/A VGND VGND VPWR VPWR _12800_/X sky130_fd_sc_hd__a2bb2o_4
X_13780_ _13779_/X VGND VGND VPWR VPWR _13780_/X sky130_fd_sc_hd__buf_2
X_22978_ _22769_/X _22974_/Y _22863_/X _22977_/X VGND VGND VPWR VPWR _22978_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_28_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12731_ _12731_/A _12731_/B VGND VGND VPWR VPWR _12731_/X sky130_fd_sc_hd__or2_4
X_24717_ _24715_/CLK _24717_/D HRESETn VGND VGND VPWR VPWR _24717_/Q sky130_fd_sc_hd__dfrtp_4
X_21929_ _21929_/A _21929_/B VGND VGND VPWR VPWR _21929_/X sky130_fd_sc_hd__or2_4
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15450_ _13899_/X _15449_/X _15446_/X _24954_/Q _15444_/X VGND VGND VPWR VPWR _24954_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_19_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12662_ _12631_/B _12659_/B _12662_/C VGND VGND VPWR VPWR _12662_/X sky130_fd_sc_hd__or3_4
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24648_ _24649_/CLK _24648_/D HRESETn VGND VGND VPWR VPWR _16230_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_128_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_101_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_203_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _20968_/A _14394_/X _14400_/X _14384_/A VGND VGND VPWR VPWR _14401_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22114__B2 _21549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15380_/X VGND VGND VPWR VPWR _15382_/B sky130_fd_sc_hd__inv_2
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12623_/A _24872_/Q _12623_/A _24872_/Q VGND VGND VPWR VPWR _12593_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22665__A2 _21413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24579_ _24572_/CLK _24579_/D HRESETn VGND VGND VPWR VPWR _22608_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24247__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ _17120_/A _17119_/X VGND VGND VPWR VPWR _17120_/X sky130_fd_sc_hd__or2_4
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _25155_/Q _14325_/X _14331_/Y VGND VGND VPWR VPWR _14332_/X sky130_fd_sc_hd__o21a_4
XFILLER_15_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_5_21_0_HCLK_A clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17051_ _17022_/Y _17051_/B VGND VGND VPWR VPWR _17053_/B sky130_fd_sc_hd__nor2_4
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _14263_/A VGND VGND VPWR VPWR _14263_/Y sky130_fd_sc_hd__inv_2
X_16002_ _15995_/X VGND VGND VPWR VPWR _16002_/X sky130_fd_sc_hd__buf_2
XFILLER_137_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13214_ _13373_/A _13214_/B VGND VGND VPWR VPWR _13215_/C sky130_fd_sc_hd__or2_4
XANTENNA__21625__B1 _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21198__A _20335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14194_ _14194_/A VGND VGND VPWR VPWR _14195_/B sky130_fd_sc_hd__buf_2
XFILLER_125_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23090__A2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13145_ _13233_/A VGND VGND VPWR VPWR _13168_/A sky130_fd_sc_hd__buf_2
XFILLER_124_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13076_ _13076_/A _13076_/B _13075_/X VGND VGND VPWR VPWR _13076_/X sky130_fd_sc_hd__and3_4
X_17953_ _17956_/A _17953_/B VGND VGND VPWR VPWR _17954_/C sky130_fd_sc_hd__or2_4
XFILLER_78_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12027_ _13527_/B _12026_/X _25293_/Q _12027_/D VGND VGND VPWR VPWR _12028_/A sky130_fd_sc_hd__or4_4
X_16904_ _16896_/X _16904_/B _16904_/C _16904_/D VGND VGND VPWR VPWR _16904_/X sky130_fd_sc_hd__or4_4
XANTENNA__25035__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17884_ _17737_/X _17878_/B _17883_/Y VGND VGND VPWR VPWR _24246_/D sky130_fd_sc_hd__and3_4
XFILLER_66_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16804__B1 HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19623_ _19621_/Y _19619_/X _19622_/X _19619_/X VGND VGND VPWR VPWR _23665_/D sky130_fd_sc_hd__a2bb2o_4
X_16835_ _16834_/Y _16830_/X _15750_/X _16830_/X VGND VGND VPWR VPWR _16835_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19554_ _19551_/Y _19552_/X _19553_/X _19552_/X VGND VGND VPWR VPWR _19554_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13978_ _13977_/X VGND VGND VPWR VPWR _13984_/A sky130_fd_sc_hd__inv_2
X_16766_ _15019_/Y _16764_/X _15747_/X _16764_/X VGND VGND VPWR VPWR _16766_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21156__A2 _15852_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18505_ _18479_/X _18496_/X _18457_/Y VGND VGND VPWR VPWR _18505_/X sky130_fd_sc_hd__o21a_4
XFILLER_19_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21661__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12929_ _12924_/A _12902_/X _12874_/X _12926_/B VGND VGND VPWR VPWR _12930_/A sky130_fd_sc_hd__a211o_4
X_15717_ _15763_/A VGND VGND VPWR VPWR _15721_/A sky130_fd_sc_hd__buf_2
X_16697_ _16697_/A VGND VGND VPWR VPWR _16697_/Y sky130_fd_sc_hd__inv_2
X_19485_ _23710_/Q VGND VGND VPWR VPWR _21483_/B sky130_fd_sc_hd__inv_2
XANTENNA__20903__A2 _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18436_ _18432_/X _18433_/X _18434_/X _18436_/D VGND VGND VPWR VPWR _18450_/B sky130_fd_sc_hd__or4_4
X_15648_ _15648_/A VGND VGND VPWR VPWR _15649_/A sky130_fd_sc_hd__buf_2
XANTENNA__24670__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15579_ _15579_/A VGND VGND VPWR VPWR _15579_/Y sky130_fd_sc_hd__inv_2
X_18367_ _18365_/A VGND VGND VPWR VPWR _18367_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21056__A1_N _21729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17318_ _17254_/C _17323_/B _17271_/X VGND VGND VPWR VPWR _17318_/Y sky130_fd_sc_hd__a21oi_4
X_18298_ _18291_/X VGND VGND VPWR VPWR _18298_/X sky130_fd_sc_hd__buf_2
XFILLER_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17249_ _24340_/Q VGND VGND VPWR VPWR _17249_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19809__B1 _19758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15543__B1 HADDR[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20260_ _20258_/Y _20254_/X _16872_/A _20259_/X VGND VGND VPWR VPWR _23434_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20191_ _20203_/A VGND VGND VPWR VPWR _20191_/X sky130_fd_sc_hd__buf_2
XANTENNA__12523__A _24852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23950_ _25098_/CLK _23950_/D HRESETn VGND VGND VPWR VPWR _23950_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18210__A _17928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22901_ _22900_/X VGND VGND VPWR VPWR _22901_/Y sky130_fd_sc_hd__inv_2
X_23881_ _23884_/CLK _23881_/D VGND VGND VPWR VPWR _19000_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22832_ _15122_/A _22832_/B VGND VGND VPWR VPWR _22832_/X sky130_fd_sc_hd__or2_4
XANTENNA__24758__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22763_ _22763_/A _22763_/B VGND VGND VPWR VPWR _22778_/B sky130_fd_sc_hd__and2_4
XANTENNA__12832__B2 _24776_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22386__B _22390_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24502_ _24502_/CLK _16623_/X HRESETn VGND VGND VPWR VPWR _16622_/A sky130_fd_sc_hd__dfrtp_4
X_21714_ _14268_/Y _21548_/B VGND VGND VPWR VPWR _21714_/Y sky130_fd_sc_hd__nor2_4
XFILLER_73_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25482_ _25284_/CLK _12030_/X HRESETn VGND VGND VPWR VPWR _11989_/A sky130_fd_sc_hd__dfrtp_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22694_ _24581_/Q _22298_/B VGND VGND VPWR VPWR _22694_/X sky130_fd_sc_hd__or2_4
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20895__A1_N _20882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24433_ _24995_/CLK _16793_/X HRESETn VGND VGND VPWR VPWR _16792_/A sky130_fd_sc_hd__dfrtp_4
X_21645_ _21645_/A VGND VGND VPWR VPWR _21645_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20107__B1 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24340__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23192__A1_N _17178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24364_ _24364_/CLK _24364_/D HRESETn VGND VGND VPWR VPWR _24364_/Q sky130_fd_sc_hd__dfrtp_4
X_21576_ _16618_/Y _21570_/X _21573_/X _21575_/X VGND VGND VPWR VPWR _21576_/X sky130_fd_sc_hd__o22a_4
XFILLER_123_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23315_ _17264_/Y _22475_/X _12859_/A _22435_/X VGND VGND VPWR VPWR _23315_/X sky130_fd_sc_hd__a2bb2o_4
X_20527_ _20428_/C _20495_/X _20443_/D _14495_/X _20433_/X VGND VGND VPWR VPWR _24078_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_138_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15534__B1 HADDR[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24295_ _25433_/CLK _17644_/X HRESETn VGND VGND VPWR VPWR _24295_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23246_ _23246_/A _21017_/B VGND VGND VPWR VPWR _23246_/X sky130_fd_sc_hd__or2_4
X_20458_ _20458_/A _20458_/B _20455_/X _20458_/D VGND VGND VPWR VPWR _24079_/D sky130_fd_sc_hd__or4_4
XFILLER_84_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12433__A _12433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23177_ _23155_/X _23158_/X _23162_/Y _23176_/X VGND VGND VPWR VPWR HRDATA[26] sky130_fd_sc_hd__a211o_4
X_20389_ _21969_/A _20386_/Y _15766_/X _20386_/Y VGND VGND VPWR VPWR _23384_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15837__A1 _15824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22128_ _15625_/A _15708_/A VGND VGND VPWR VPWR _22128_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_26_0_HCLK clkbuf_7_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_14950_ _14949_/Y _24415_/Q _14949_/Y _24415_/Q VGND VGND VPWR VPWR _14950_/X sky130_fd_sc_hd__a2bb2o_4
X_22059_ _22050_/X _19270_/Y VGND VGND VPWR VPWR _22059_/X sky130_fd_sc_hd__or2_4
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_89_0_HCLK clkbuf_6_44_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_89_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13901_ _24952_/Q VGND VGND VPWR VPWR _13901_/X sky130_fd_sc_hd__buf_2
X_14881_ _14881_/A VGND VGND VPWR VPWR _14881_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13832_ _13831_/Y _13829_/X _11825_/X _13829_/X VGND VGND VPWR VPWR _25251_/D sky130_fd_sc_hd__a2bb2o_4
X_16620_ _16620_/A VGND VGND VPWR VPWR _16620_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16586__A1_N _16585_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24499__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16551_ _16558_/A VGND VGND VPWR VPWR _16551_/X sky130_fd_sc_hd__buf_2
XFILLER_95_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13763_ _13763_/A VGND VGND VPWR VPWR _14703_/A sky130_fd_sc_hd__buf_2
XFILLER_95_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22886__A2 _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24428__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ _12708_/A _12708_/B VGND VGND VPWR VPWR _12714_/Y sky130_fd_sc_hd__nand2_4
X_15502_ _15501_/Y _15499_/X HADDR[18] _15499_/X VGND VGND VPWR VPWR _24930_/D sky130_fd_sc_hd__a2bb2o_4
X_16482_ _16481_/Y _16479_/X _16306_/X _16479_/X VGND VGND VPWR VPWR _16482_/X sky130_fd_sc_hd__a2bb2o_4
X_19270_ _23786_/Q VGND VGND VPWR VPWR _19270_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13694_ _13693_/X _13694_/B VGND VGND VPWR VPWR _13695_/B sky130_fd_sc_hd__or2_4
XFILLER_43_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15433_ _15430_/X VGND VGND VPWR VPWR _15452_/A sky130_fd_sc_hd__inv_2
X_18221_ _18221_/A _19193_/A VGND VGND VPWR VPWR _18223_/B sky130_fd_sc_hd__or2_4
XFILLER_54_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12645_ _12645_/A _12645_/B VGND VGND VPWR VPWR _12645_/X sky130_fd_sc_hd__or2_4
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16725__D _21314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24081__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ _15296_/A _15362_/X _15363_/Y VGND VGND VPWR VPWR _24982_/D sky130_fd_sc_hd__o21a_4
X_18152_ _18184_/A _18150_/X _18152_/C VGND VGND VPWR VPWR _18153_/C sky130_fd_sc_hd__and3_4
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12576_ _25403_/Q VGND VGND VPWR VPWR _12576_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24010__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14315_ _25162_/Q _14302_/X _25161_/Q _14307_/X VGND VGND VPWR VPWR _14315_/X sky130_fd_sc_hd__o22a_4
X_17103_ _16972_/Y _17108_/B _17056_/X VGND VGND VPWR VPWR _17103_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18083_ _18221_/A _18083_/B VGND VGND VPWR VPWR _18083_/X sky130_fd_sc_hd__or2_4
XANTENNA__15525__B1 HADDR[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15295_ _24984_/Q VGND VGND VPWR VPWR _15356_/A sky130_fd_sc_hd__inv_2
X_17034_ _17034_/A _17034_/B _17033_/X VGND VGND VPWR VPWR _17034_/X sky130_fd_sc_hd__or3_4
X_14246_ _13964_/X _14245_/X VGND VGND VPWR VPWR _15441_/A sky130_fd_sc_hd__or2_4
XFILLER_7_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23063__A2 _22998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25287__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14177_ _25118_/Q VGND VGND VPWR VPWR _14177_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25216__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13128_ _13128_/A _13128_/B VGND VGND VPWR VPWR _13129_/B sky130_fd_sc_hd__or2_4
XFILLER_113_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18985_ _18984_/Y _18972_/A _17443_/X _18972_/A VGND VGND VPWR VPWR _23885_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13059_ _13054_/A _13062_/B VGND VGND VPWR VPWR _13059_/Y sky130_fd_sc_hd__nand2_4
X_17936_ _17931_/X _17935_/X _18017_/A VGND VGND VPWR VPWR _17944_/B sky130_fd_sc_hd__o21a_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17867_ _17867_/A _17867_/B VGND VGND VPWR VPWR _17867_/X sky130_fd_sc_hd__or2_4
XFILLER_94_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15056__A2 _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17176__A2_N _17350_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19606_ _23669_/Q VGND VGND VPWR VPWR _19606_/Y sky130_fd_sc_hd__inv_2
X_16818_ _14969_/Y _16816_/X HWDATA[20] _16816_/X VGND VGND VPWR VPWR _16818_/X sky130_fd_sc_hd__a2bb2o_4
X_17798_ _17738_/X _17796_/X _17798_/C VGND VGND VPWR VPWR _17798_/X sky130_fd_sc_hd__and3_4
XANTENNA__24851__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19537_ _16725_/A _16725_/B _13775_/X _19536_/Y VGND VGND VPWR VPWR _19538_/A sky130_fd_sc_hd__and4_4
X_16749_ _16739_/A VGND VGND VPWR VPWR _16749_/X sky130_fd_sc_hd__buf_2
XANTENNA__16485__A _16485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12814__B2 _24787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19468_ _17708_/A _17713_/A _19492_/B VGND VGND VPWR VPWR _19888_/C sky130_fd_sc_hd__or3_4
XANTENNA__18950__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18419_ _24636_/Q _24147_/Q _16263_/Y _18418_/Y VGND VGND VPWR VPWR _18419_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15764__B1 _15627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19399_ _14656_/Y _19038_/B _19399_/C VGND VGND VPWR VPWR _19400_/A sky130_fd_sc_hd__or3_4
XFILLER_37_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21430_ _21062_/Y VGND VGND VPWR VPWR _22963_/A sky130_fd_sc_hd__buf_2
XFILLER_33_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21361_ _21332_/Y _21343_/X _21349_/Y _21360_/Y VGND VGND VPWR VPWR _21361_/X sky130_fd_sc_hd__a211o_4
X_23100_ _23100_/A VGND VGND VPWR VPWR _23274_/A sky130_fd_sc_hd__buf_2
X_20312_ _20310_/Y _20311_/X _19992_/X _20311_/X VGND VGND VPWR VPWR _20312_/X sky130_fd_sc_hd__a2bb2o_4
X_24080_ _23995_/CLK _24080_/D HRESETn VGND VGND VPWR VPWR _20426_/B sky130_fd_sc_hd__dfrtp_4
X_21292_ _21071_/A VGND VGND VPWR VPWR _21293_/A sky130_fd_sc_hd__buf_2
X_23031_ _24758_/Q _23140_/B VGND VGND VPWR VPWR _23031_/X sky130_fd_sc_hd__or2_4
X_20243_ _20242_/Y _20238_/X _19740_/X _20238_/X VGND VGND VPWR VPWR _23440_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22262__B1 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20174_ _20174_/A VGND VGND VPWR VPWR _20174_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24982_ _24980_/CLK _24982_/D HRESETn VGND VGND VPWR VPWR _24982_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23933_ _23933_/CLK _23933_/D HRESETn VGND VGND VPWR VPWR _23933_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23864_ _25485_/CLK _23864_/D VGND VGND VPWR VPWR _19049_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24592__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22815_ _22815_/A _21048_/B VGND VGND VPWR VPWR _22815_/X sky130_fd_sc_hd__or2_4
XANTENNA__20328__B1 _15766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23795_ _24398_/CLK _23795_/D VGND VGND VPWR VPWR _19246_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__19194__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24521__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25534_ _24691_/CLK _11758_/X HRESETn VGND VGND VPWR VPWR _11756_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_38_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23005__B _22810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22746_ _22544_/X _22745_/X _22466_/A _25522_/Q _22922_/A VGND VGND VPWR VPWR _22746_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18613__A1_N _24523_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18941__B1 _18940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15755__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25465_ _24368_/CLK _12103_/X HRESETn VGND VGND VPWR VPWR _12092_/A sky130_fd_sc_hd__dfrtp_4
X_22677_ _16687_/Y _22677_/B VGND VGND VPWR VPWR _22677_/X sky130_fd_sc_hd__and2_4
XFILLER_41_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12430_ _12430_/A _12235_/X _12283_/X _12382_/X VGND VGND VPWR VPWR _12430_/X sky130_fd_sc_hd__or4_4
X_24416_ _24462_/CLK _16828_/X HRESETn VGND VGND VPWR VPWR _24416_/Q sky130_fd_sc_hd__dfrtp_4
X_21628_ _21609_/A _21628_/B _21628_/C VGND VGND VPWR VPWR _21628_/X sky130_fd_sc_hd__and3_4
X_25396_ _25397_/CLK _12717_/X HRESETn VGND VGND VPWR VPWR _25396_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23293__A2 _22467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23021__A _23021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12361_ _25344_/Q VGND VGND VPWR VPWR _12999_/B sky130_fd_sc_hd__inv_2
XFILLER_138_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15739__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15507__B1 HADDR[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24347_ _24345_/CLK _17319_/X HRESETn VGND VGND VPWR VPWR _17192_/A sky130_fd_sc_hd__dfrtp_4
X_21559_ _21559_/A _13467_/X VGND VGND VPWR VPWR _21559_/X sky130_fd_sc_hd__or2_4
XFILLER_138_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14100_ _14100_/A _14100_/B _14115_/A VGND VGND VPWR VPWR _14101_/B sky130_fd_sc_hd__or3_4
X_15080_ _15080_/A VGND VGND VPWR VPWR _15080_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16338__A2_N _16337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12292_ _25333_/Q VGND VGND VPWR VPWR _12292_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25380__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24278_ _24278_/CLK _17699_/Y HRESETn VGND VGND VPWR VPWR _17577_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14031_ _14031_/A VGND VGND VPWR VPWR _14070_/B sky130_fd_sc_hd__inv_2
XANTENNA__21056__B2 _21729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23229_ _23124_/A _23229_/B VGND VGND VPWR VPWR _23229_/Y sky130_fd_sc_hd__nor2_4
XFILLER_10_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21476__A _21454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15474__A _16359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18770_ _18765_/A _18765_/B _18733_/X _18767_/B VGND VGND VPWR VPWR _18771_/A sky130_fd_sc_hd__a211o_4
X_15982_ _15937_/Y VGND VGND VPWR VPWR _15982_/X sky130_fd_sc_hd__buf_2
XFILLER_122_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17721_ _17720_/X VGND VGND VPWR VPWR _17722_/A sky130_fd_sc_hd__buf_2
XFILLER_0_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14933_ _15063_/A VGND VGND VPWR VPWR _15262_/A sky130_fd_sc_hd__buf_2
XFILLER_76_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24609__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17652_ _17624_/A VGND VGND VPWR VPWR _17652_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_113_0_HCLK clkbuf_7_56_0_HCLK/X VGND VGND VPWR VPWR _24541_/CLK sky130_fd_sc_hd__clkbuf_1
X_14864_ _14869_/A _14798_/B _14870_/A _14880_/B VGND VGND VPWR VPWR _14864_/X sky130_fd_sc_hd__or4_4
XFILLER_75_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16603_ _16603_/A VGND VGND VPWR VPWR _16603_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_176_0_HCLK clkbuf_7_88_0_HCLK/X VGND VGND VPWR VPWR _24288_/CLK sky130_fd_sc_hd__clkbuf_1
X_13815_ _13815_/A _17413_/A VGND VGND VPWR VPWR _13815_/X sky130_fd_sc_hd__or2_4
X_14795_ _20995_/B VGND VGND VPWR VPWR _20996_/B sky130_fd_sc_hd__inv_2
X_17583_ _17560_/Y _17582_/X VGND VGND VPWR VPWR _17583_/X sky130_fd_sc_hd__or2_4
XFILLER_21_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24262__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19322_ _23768_/Q VGND VGND VPWR VPWR _19322_/Y sky130_fd_sc_hd__inv_2
X_13746_ _13746_/A VGND VGND VPWR VPWR _13763_/A sky130_fd_sc_hd__inv_2
X_16534_ _16533_/Y _16531_/X _16359_/X _16531_/X VGND VGND VPWR VPWR _24537_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19253_ _23792_/Q VGND VGND VPWR VPWR _19253_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16455__D _21314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13677_ _13695_/A VGND VGND VPWR VPWR _13713_/A sky130_fd_sc_hd__inv_2
X_16465_ _24563_/Q VGND VGND VPWR VPWR _16465_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15746__B1 _24856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18204_ _18204_/A _18204_/B VGND VGND VPWR VPWR _18205_/C sky130_fd_sc_hd__or2_4
X_12628_ _12664_/A VGND VGND VPWR VPWR _12631_/B sky130_fd_sc_hd__inv_2
X_15416_ _15159_/X _15415_/X VGND VGND VPWR VPWR _15416_/Y sky130_fd_sc_hd__nand2_4
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16396_ _24590_/Q VGND VGND VPWR VPWR _16396_/Y sky130_fd_sc_hd__inv_2
X_19184_ _19183_/Y _19181_/X _19071_/X _19181_/X VGND VGND VPWR VPWR _23817_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25468__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15347_ _15306_/X _15316_/X _15336_/C VGND VGND VPWR VPWR _15347_/X sky130_fd_sc_hd__o21a_4
X_18135_ _18066_/A _23767_/Q VGND VGND VPWR VPWR _18135_/X sky130_fd_sc_hd__or2_4
X_12559_ _12559_/A VGND VGND VPWR VPWR _12559_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14553__A HREADY VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15278_ _15278_/A _15278_/B VGND VGND VPWR VPWR _15282_/B sky130_fd_sc_hd__or2_4
X_18066_ _18066_/A _18066_/B VGND VGND VPWR VPWR _18068_/B sky130_fd_sc_hd__or2_4
XFILLER_32_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22770__A _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14229_ _14224_/A VGND VGND VPWR VPWR _14229_/X sky130_fd_sc_hd__buf_2
X_17017_ _16998_/X _17003_/X _17017_/C _17017_/D VGND VGND VPWR VPWR _17017_/X sky130_fd_sc_hd__or4_4
XANTENNA__25050__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12073__A _12072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18999__B1 _18997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18968_ _18967_/Y _14665_/X _17418_/X _14665_/X VGND VGND VPWR VPWR _18968_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12801__A _22706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17919_ _13541_/B VGND VGND VPWR VPWR _17920_/B sky130_fd_sc_hd__inv_2
X_18899_ _13755_/A _13748_/A _13746_/A VGND VGND VPWR VPWR _19822_/C sky130_fd_sc_hd__or3_4
Xclkbuf_7_72_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_72_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20930_ _20931_/B VGND VGND VPWR VPWR _20930_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14237__B1 _13803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23106__A _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20861_ _13661_/B VGND VGND VPWR VPWR _20861_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15985__B1 _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22600_ _21580_/A _22600_/B VGND VGND VPWR VPWR _22600_/Y sky130_fd_sc_hd__nor2_4
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23580_ _23580_/CLK _19869_/X VGND VGND VPWR VPWR _19865_/A sky130_fd_sc_hd__dfxtp_4
X_20792_ _20790_/A _20787_/X VGND VGND VPWR VPWR _20792_/X sky130_fd_sc_hd__or2_4
XFILLER_126_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22531_ _13580_/Y _22531_/B VGND VGND VPWR VPWR _22531_/X sky130_fd_sc_hd__and2_4
XFILLER_39_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15737__B1 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22664__B _22664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23985__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25250_ _25263_/CLK _13834_/X HRESETn VGND VGND VPWR VPWR _13575_/A sky130_fd_sc_hd__dfrtp_4
X_22462_ _22462_/A _22462_/B _22462_/C _22462_/D VGND VGND VPWR VPWR _22462_/X sky130_fd_sc_hd__or4_4
XFILLER_37_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17758__B _17758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24201_ _24290_/CLK _18302_/X HRESETn VGND VGND VPWR VPWR _24201_/Q sky130_fd_sc_hd__dfrtp_4
X_21413_ _23034_/A VGND VGND VPWR VPWR _21413_/X sky130_fd_sc_hd__buf_2
XANTENNA__22383__C _22383_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25181_ _24148_/CLK _14242_/X HRESETn VGND VGND VPWR VPWR _25181_/Q sky130_fd_sc_hd__dfstp_4
X_22393_ _22523_/A VGND VGND VPWR VPWR _22393_/X sky130_fd_sc_hd__buf_2
XANTENNA__25138__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24132_ _24555_/CLK _24132_/D HRESETn VGND VGND VPWR VPWR _24132_/Q sky130_fd_sc_hd__dfrtp_4
X_21344_ SSn_S3 _12054_/X SSn_S2 _13468_/X VGND VGND VPWR VPWR _21344_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16162__B1 _15986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24063_ _25397_/CLK _24063_/D HRESETn VGND VGND VPWR VPWR _15484_/A sky130_fd_sc_hd__dfrtp_4
X_21275_ _21103_/X VGND VGND VPWR VPWR _21275_/X sky130_fd_sc_hd__buf_2
XFILLER_85_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12414__C _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23014_ _24051_/Q _21287_/Y _24019_/Q _21589_/X VGND VGND VPWR VPWR _23014_/Y sky130_fd_sc_hd__a22oi_4
X_20226_ _20226_/A VGND VGND VPWR VPWR _20226_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20157_ _20156_/Y _20154_/X _20089_/X _20154_/X VGND VGND VPWR VPWR _20157_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24773__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24965_ _24977_/CLK _24965_/D HRESETn VGND VGND VPWR VPWR _15114_/A sky130_fd_sc_hd__dfrtp_4
X_20088_ _23497_/Q VGND VGND VPWR VPWR _20088_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12430__B _12235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24702__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11930_ _19612_/A VGND VGND VPWR VPWR _11930_/X sky130_fd_sc_hd__buf_2
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23916_ _24398_/CLK _18903_/X VGND VGND VPWR VPWR _18897_/A sky130_fd_sc_hd__dfxtp_4
X_24896_ _24018_/CLK _15598_/X HRESETn VGND VGND VPWR VPWR _15597_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11861_ HWDATA[1] VGND VGND VPWR VPWR _11862_/A sky130_fd_sc_hd__buf_2
X_23847_ _23847_/CLK _19099_/X VGND VGND VPWR VPWR _23847_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15976__B1 _15897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_249_0_HCLK clkbuf_7_124_0_HCLK/X VGND VGND VPWR VPWR _24847_/CLK sky130_fd_sc_hd__clkbuf_1
X_13600_ _14659_/A VGND VGND VPWR VPWR _19038_/D sky130_fd_sc_hd__inv_2
XFILLER_14_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14580_ _14582_/B VGND VGND VPWR VPWR _14581_/B sky130_fd_sc_hd__inv_2
X_11792_ _11790_/Y _11785_/X _11791_/X _11785_/X VGND VGND VPWR VPWR _25524_/D sky130_fd_sc_hd__a2bb2o_4
X_23778_ _23618_/CLK _19296_/X VGND VGND VPWR VPWR _13282_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_53_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12591__A2_N _24845_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13531_ _20955_/B _13530_/X SCLK_S2 _20955_/B VGND VGND VPWR VPWR _25292_/D sky130_fd_sc_hd__a2bb2o_4
X_25517_ _24285_/CLK _11823_/X HRESETn VGND VGND VPWR VPWR _25517_/Q sky130_fd_sc_hd__dfrtp_4
X_22729_ _24044_/Q _21302_/A _24012_/Q _21304_/X VGND VGND VPWR VPWR _22729_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16250_ _16249_/Y _16247_/X _16147_/X _16247_/X VGND VGND VPWR VPWR _24642_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13462_ _13177_/Y _13454_/X _13461_/X VGND VGND VPWR VPWR _13462_/X sky130_fd_sc_hd__and3_4
X_25448_ _25449_/CLK _25448_/D HRESETn VGND VGND VPWR VPWR _25448_/Q sky130_fd_sc_hd__dfrtp_4
X_15201_ _15201_/A VGND VGND VPWR VPWR _15201_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12413_ _12413_/A VGND VGND VPWR VPWR _12413_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16181_ _16180_/X VGND VGND VPWR VPWR _16449_/A sky130_fd_sc_hd__buf_2
X_13393_ _13457_/A _13393_/B _13392_/X VGND VGND VPWR VPWR _13397_/B sky130_fd_sc_hd__and3_4
X_25379_ _25385_/CLK _25379_/D HRESETn VGND VGND VPWR VPWR _12771_/A sky130_fd_sc_hd__dfrtp_4
X_15132_ _15124_/X _15127_/X _15129_/X _15131_/X VGND VGND VPWR VPWR _15132_/X sky130_fd_sc_hd__or4_4
X_12344_ _24808_/Q VGND VGND VPWR VPWR _12344_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16153__B1 _16061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22590__A _24746_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15063_ _15063_/A _15063_/B _15251_/C _15248_/A VGND VGND VPWR VPWR _15063_/X sky130_fd_sc_hd__or4_4
X_19940_ _23552_/Q VGND VGND VPWR VPWR _21796_/B sky130_fd_sc_hd__inv_2
X_12275_ _12509_/A VGND VGND VPWR VPWR _12389_/A sky130_fd_sc_hd__buf_2
XFILLER_5_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14014_ _14010_/X _14013_/Y _14010_/X _14013_/Y VGND VGND VPWR VPWR _14538_/D sky130_fd_sc_hd__a2bb2o_4
X_19871_ _19870_/Y _19868_/X _19615_/X _19868_/X VGND VGND VPWR VPWR _19871_/X sky130_fd_sc_hd__a2bb2o_4
X_18822_ _18742_/A _18783_/X _18822_/C VGND VGND VPWR VPWR _24113_/D sky130_fd_sc_hd__and3_4
XANTENNA__16456__B2 _16455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14204__A1_N _20500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18753_ _18758_/A _18757_/A _18753_/C _18756_/B VGND VGND VPWR VPWR _18759_/B sky130_fd_sc_hd__or4_4
XFILLER_110_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21934__A _21455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15965_ _12228_/Y _15960_/X _15964_/X _15960_/X VGND VGND VPWR VPWR _15965_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11882__D _13678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24443__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17704_ _24200_/Q VGND VGND VPWR VPWR _21194_/A sky130_fd_sc_hd__buf_2
XFILLER_49_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_59_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14916_ _24409_/Q VGND VGND VPWR VPWR _14916_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19404__A _19642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18684_ _18623_/Y _18782_/A _18680_/X _18683_/X VGND VGND VPWR VPWR _18693_/A sky130_fd_sc_hd__or4_4
X_15896_ _15900_/A VGND VGND VPWR VPWR _15896_/X sky130_fd_sc_hd__buf_2
X_17635_ _17565_/Y _17635_/B VGND VGND VPWR VPWR _17645_/B sky130_fd_sc_hd__or2_4
X_14847_ _14846_/X VGND VGND VPWR VPWR _14847_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19158__B1 _19133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17566_ _24292_/Q VGND VGND VPWR VPWR _17567_/D sky130_fd_sc_hd__inv_2
X_14778_ _14778_/A VGND VGND VPWR VPWR _14778_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19305_ _19304_/Y _19302_/X _19191_/X _19302_/X VGND VGND VPWR VPWR _19305_/X sky130_fd_sc_hd__a2bb2o_4
X_16517_ _16515_/Y _16511_/X _16143_/X _16516_/X VGND VGND VPWR VPWR _24543_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13729_ _13729_/A _13729_/B VGND VGND VPWR VPWR _13729_/Y sky130_fd_sc_hd__nand2_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15719__B1 _11749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17859__A _17846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17497_ _17497_/A _17497_/B _17495_/X _17497_/D VGND VGND VPWR VPWR _17497_/X sky130_fd_sc_hd__or4_4
XANTENNA__16763__A _24447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22484__B _22644_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19236_ _19234_/Y _19235_/X _19212_/X _19235_/X VGND VGND VPWR VPWR _19236_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16448_ _16448_/A VGND VGND VPWR VPWR _18496_/A sky130_fd_sc_hd__buf_2
XANTENNA__16392__B1 _16300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23299__C _23299_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15379__A _15336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19167_ _19153_/Y VGND VGND VPWR VPWR _19167_/X sky130_fd_sc_hd__buf_2
XFILLER_118_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16913__D _16913_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16379_ _16378_/Y _16375_/X _16285_/X _16375_/X VGND VGND VPWR VPWR _24597_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25231__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19330__B1 _19307_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18118_ _18221_/A _18118_/B VGND VGND VPWR VPWR _18118_/X sky130_fd_sc_hd__or2_4
XFILLER_69_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19098_ _19098_/A VGND VGND VPWR VPWR _19098_/X sky130_fd_sc_hd__buf_2
XFILLER_117_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18049_ _18177_/A VGND VGND VPWR VPWR _18058_/A sky130_fd_sc_hd__buf_2
X_21060_ _11864_/A _21049_/X _21050_/X _21059_/X VGND VGND VPWR VPWR _21060_/X sky130_fd_sc_hd__a211o_4
XFILLER_63_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20011_ _23528_/Q VGND VGND VPWR VPWR _21793_/B sky130_fd_sc_hd__inv_2
XFILLER_115_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21728__C1 _21727_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24184__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19397__B1 _19307_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22659__B _22534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24750_ _24766_/CLK _24750_/D HRESETn VGND VGND VPWR VPWR _24750_/Q sky130_fd_sc_hd__dfrtp_4
X_21962_ _21962_/A _19598_/A VGND VGND VPWR VPWR _21962_/X sky130_fd_sc_hd__and2_4
XFILLER_55_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24113__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23701_ _23396_/CLK _19512_/X VGND VGND VPWR VPWR _19511_/A sky130_fd_sc_hd__dfxtp_4
X_20913_ _20913_/A VGND VGND VPWR VPWR _20913_/X sky130_fd_sc_hd__buf_2
XANTENNA__15958__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24681_ _24682_/CLK _24681_/D HRESETn VGND VGND VPWR VPWR _22655_/A sky130_fd_sc_hd__dfrtp_4
X_21893_ _21890_/X _21891_/X _21893_/C VGND VGND VPWR VPWR _21893_/X sky130_fd_sc_hd__and3_4
XFILLER_55_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20951__B1 _11958_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23632_ _23649_/CLK _23632_/D VGND VGND VPWR VPWR _19717_/A sky130_fd_sc_hd__dfxtp_4
X_20844_ _20843_/X VGND VGND VPWR VPWR _24035_/D sky130_fd_sc_hd__inv_2
XFILLER_42_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_2_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15973__A3 _11812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_16_0_HCLK clkbuf_7_8_0_HCLK/X VGND VGND VPWR VPWR _25309_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23563_ _23516_/CLK _19914_/X VGND VGND VPWR VPWR _23563_/Q sky130_fd_sc_hd__dfxtp_4
X_20775_ _20770_/X _20773_/X _24901_/Q _20774_/X VGND VGND VPWR VPWR _20775_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25319__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_79_0_HCLK clkbuf_8_79_0_HCLK/A VGND VGND VPWR VPWR _24148_/CLK sky130_fd_sc_hd__clkbuf_1
X_25302_ _25290_/CLK _25302_/D HRESETn VGND VGND VPWR VPWR _12014_/A sky130_fd_sc_hd__dfrtp_4
X_22514_ _22278_/X _22512_/X _21106_/X _22513_/X VGND VGND VPWR VPWR _22514_/X sky130_fd_sc_hd__o22a_4
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16383__B1 _16380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23248__A2 _21021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23494_ _23494_/CLK _20100_/X VGND VGND VPWR VPWR _23494_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25233_ _24643_/CLK _13879_/X HRESETn VGND VGND VPWR VPWR _25233_/Q sky130_fd_sc_hd__dfrtp_4
X_22445_ _16518_/Y _21067_/X _16728_/A _16603_/Y _16795_/A VGND VGND VPWR VPWR _22445_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__23002__C _23002_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19321__B1 _19206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11747__B2 _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25164_ _25309_/CLK _25164_/D HRESETn VGND VGND VPWR VPWR _25164_/Q sky130_fd_sc_hd__dfrtp_4
X_22376_ _22068_/A _22376_/B VGND VGND VPWR VPWR _22376_/X sky130_fd_sc_hd__or2_4
XFILLER_124_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24115_ _24120_/CLK _24115_/D HRESETn VGND VGND VPWR VPWR _18633_/A sky130_fd_sc_hd__dfrtp_4
X_21327_ _24535_/Q _22592_/B _21326_/X VGND VGND VPWR VPWR _21327_/X sky130_fd_sc_hd__o21a_4
XFILLER_89_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20482__A2 _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21738__B _21582_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25095_ _25137_/CLK _14520_/X HRESETn VGND VGND VPWR VPWR _25095_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24954__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12060_ _13533_/A _12060_/B _15652_/D _12059_/X VGND VGND VPWR VPWR _12060_/X sky130_fd_sc_hd__or4_4
X_24046_ _24049_/CLK _20895_/X HRESETn VGND VGND VPWR VPWR _24046_/Q sky130_fd_sc_hd__dfrtp_4
X_21258_ _21254_/X _21257_/X _14676_/X VGND VGND VPWR VPWR _21259_/C sky130_fd_sc_hd__o21a_4
XFILLER_2_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20209_ _20209_/A VGND VGND VPWR VPWR _20209_/Y sky130_fd_sc_hd__inv_2
X_21189_ _21184_/A _20356_/Y VGND VGND VPWR VPWR _21191_/B sky130_fd_sc_hd__or2_4
XFILLER_77_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21982__A2 _21911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15752__A HWDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12962_ _12774_/Y _12964_/B _12961_/Y VGND VGND VPWR VPWR _12962_/X sky130_fd_sc_hd__o21a_4
X_15750_ HWDATA[12] VGND VGND VPWR VPWR _15750_/X sky130_fd_sc_hd__buf_2
X_24948_ _24950_/CLK _24948_/D HRESETn VGND VGND VPWR VPWR _13927_/D sky130_fd_sc_hd__dfrtp_4
X_11913_ _11870_/A _11884_/X _11916_/B _11878_/A _11912_/Y VGND VGND VPWR VPWR _11913_/X
+ sky130_fd_sc_hd__a32o_4
X_14701_ _20043_/A _14684_/A _13735_/X _14746_/A VGND VGND VPWR VPWR _14701_/X sky130_fd_sc_hd__o22a_4
XFILLER_73_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12893_ _12841_/B _12887_/X _12874_/X _12890_/B VGND VGND VPWR VPWR _12894_/A sky130_fd_sc_hd__a211o_4
X_15681_ _15681_/A VGND VGND VPWR VPWR _15687_/B sky130_fd_sc_hd__inv_2
X_24879_ _24026_/CLK _24879_/D HRESETn VGND VGND VPWR VPWR _21008_/B sky130_fd_sc_hd__dfrtp_4
X_17420_ _17420_/A VGND VGND VPWR VPWR _17420_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13272__A _13310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11844_ _25511_/Q VGND VGND VPWR VPWR _11844_/Y sky130_fd_sc_hd__inv_2
X_14632_ _14632_/A _14616_/X VGND VGND VPWR VPWR _14632_/X sky130_fd_sc_hd__or2_4
XFILLER_61_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14563_ _13582_/Y _14563_/B VGND VGND VPWR VPWR _14601_/B sky130_fd_sc_hd__or2_4
X_17351_ _17353_/B VGND VGND VPWR VPWR _17352_/B sky130_fd_sc_hd__inv_2
X_11775_ _11773_/Y _11768_/X _11774_/X _11768_/X VGND VGND VPWR VPWR _11775_/X sky130_fd_sc_hd__a2bb2o_4
X_16302_ _23073_/A VGND VGND VPWR VPWR _16302_/Y sky130_fd_sc_hd__inv_2
X_13514_ _13514_/A VGND VGND VPWR VPWR _13514_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14494_ _13976_/X VGND VGND VPWR VPWR _14541_/A sky130_fd_sc_hd__buf_2
X_17282_ _17260_/A _17282_/B VGND VGND VPWR VPWR _17283_/A sky130_fd_sc_hd__or2_4
XFILLER_13_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19021_ _19020_/Y _19016_/X _18993_/X _19016_/X VGND VGND VPWR VPWR _23875_/D sky130_fd_sc_hd__a2bb2o_4
X_13445_ _13413_/A _13443_/X _13445_/C VGND VGND VPWR VPWR _13446_/C sky130_fd_sc_hd__and3_4
X_16233_ _16230_/Y _16225_/X _16231_/X _16232_/X VGND VGND VPWR VPWR _24648_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13376_ _13269_/A _13376_/B VGND VGND VPWR VPWR _13378_/B sky130_fd_sc_hd__or2_4
X_16164_ _16163_/Y _16088_/A _15840_/X _16088_/A VGND VGND VPWR VPWR _24669_/D sky130_fd_sc_hd__a2bb2o_4
X_12327_ _25351_/Q VGND VGND VPWR VPWR _13001_/C sky130_fd_sc_hd__inv_2
X_15115_ _15115_/A VGND VGND VPWR VPWR _15115_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16095_ _16092_/Y _16088_/X _15940_/X _16094_/X VGND VGND VPWR VPWR _16095_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15927__A _15845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18303__A _21465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24695__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15046_ _14903_/X _15025_/Y _25022_/Q _15015_/Y VGND VGND VPWR VPWR _15047_/D sky130_fd_sc_hd__a2bb2o_4
X_19923_ _19923_/A VGND VGND VPWR VPWR _19923_/X sky130_fd_sc_hd__buf_2
X_12258_ _12290_/A _24761_/Q _12260_/A _12257_/Y VGND VGND VPWR VPWR _12258_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24624__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19854_ _19854_/A VGND VGND VPWR VPWR _21899_/B sky130_fd_sc_hd__inv_2
XFILLER_116_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12189_ _12440_/C _24751_/Q _12188_/A _24751_/Q VGND VGND VPWR VPWR _12198_/A sky130_fd_sc_hd__a2bb2o_4
X_18805_ _18623_/Y _18803_/X _18804_/Y VGND VGND VPWR VPWR _18805_/X sky130_fd_sc_hd__o21a_4
X_19785_ _19782_/Y _19776_/X _19783_/X _19784_/X VGND VGND VPWR VPWR _23610_/D sky130_fd_sc_hd__a2bb2o_4
X_16997_ _16039_/Y _24374_/Q _16039_/Y _24374_/Q VGND VGND VPWR VPWR _16997_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16758__A _16733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18736_ _18736_/A VGND VGND VPWR VPWR _18737_/B sky130_fd_sc_hd__inv_2
XFILLER_62_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15948_ _15930_/X _15935_/X HWDATA[25] _24760_/Q _15933_/X VGND VGND VPWR VPWR _15948_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_95_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25121__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18667_ _18645_/X _18667_/B _18667_/C _18666_/X VGND VGND VPWR VPWR _18667_/X sky130_fd_sc_hd__or4_4
X_15879_ _15868_/X VGND VGND VPWR VPWR _15879_/X sky130_fd_sc_hd__buf_2
XANTENNA__25184__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17618_ _17618_/A VGND VGND VPWR VPWR _17618_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18598_ _16594_/Y _18789_/A _16594_/Y _18789_/A VGND VGND VPWR VPWR _18598_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25483__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22495__A _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_232_0_HCLK clkbuf_8_233_0_HCLK/A VGND VGND VPWR VPWR _25385_/CLK sky130_fd_sc_hd__clkbuf_1
X_17549_ _11835_/Y _17494_/A _11850_/Y _17573_/A VGND VGND VPWR VPWR _17549_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17589__A _17624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25412__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20560_ _20560_/A VGND VGND VPWR VPWR _23936_/D sky130_fd_sc_hd__inv_2
XFILLER_123_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19219_ _17465_/X _24194_/Q _19219_/C VGND VGND VPWR VPWR _19219_/X sky130_fd_sc_hd__or3_4
XANTENNA__22438__B1 _12202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20491_ _20491_/A _20490_/Y VGND VGND VPWR VPWR _24074_/D sky130_fd_sc_hd__or2_4
XFILLER_20_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19303__B1 _19212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22230_ _18307_/X VGND VGND VPWR VPWR _22246_/A sky130_fd_sc_hd__buf_2
XANTENNA__22989__B2 _21211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22161_ _22161_/A VGND VGND VPWR VPWR _22161_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19309__A _19309_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21112_ _21007_/A _21112_/B VGND VGND VPWR VPWR _21112_/Y sky130_fd_sc_hd__nor2_4
X_22092_ _16611_/A _21858_/X _22090_/X _22091_/X VGND VGND VPWR VPWR _22093_/C sky130_fd_sc_hd__a211o_4
XFILLER_87_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24365__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21043_ _11720_/B VGND VGND VPWR VPWR _21043_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24323__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21574__A _15852_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18290__B1 _17700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24802_ _24832_/CLK _24802_/D HRESETn VGND VGND VPWR VPWR _24802_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22994_ _24523_/Q _22922_/X _22923_/X _22993_/X VGND VGND VPWR VPWR _22995_/C sky130_fd_sc_hd__a211o_4
XFILLER_55_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_42_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_85_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21945_ _21945_/A _19621_/Y VGND VGND VPWR VPWR _21945_/X sky130_fd_sc_hd__or2_4
X_24733_ _24356_/CLK _24733_/D HRESETn VGND VGND VPWR VPWR _24733_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24664_ _24654_/CLK _16190_/X HRESETn VGND VGND VPWR VPWR _23291_/A sky130_fd_sc_hd__dfrtp_4
X_21876_ _14689_/A _19831_/Y VGND VGND VPWR VPWR _21879_/B sky130_fd_sc_hd__or2_4
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23615_ _23623_/CLK _19767_/X VGND VGND VPWR VPWR _23615_/Q sky130_fd_sc_hd__dfxtp_4
X_20827_ _20827_/A VGND VGND VPWR VPWR _20827_/Y sky130_fd_sc_hd__inv_2
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24595_ _24596_/CLK _16385_/X HRESETn VGND VGND VPWR VPWR _24595_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19542__B1 _19404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23546_ _23545_/CLK _23546_/D VGND VGND VPWR VPWR _23546_/Q sky130_fd_sc_hd__dfxtp_4
X_20758_ _13119_/A _13119_/B _13119_/C _20772_/C VGND VGND VPWR VPWR _20758_/X sky130_fd_sc_hd__or4_4
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23477_ _23494_/CLK _20145_/X VGND VGND VPWR VPWR _20144_/A sky130_fd_sc_hd__dfxtp_4
X_20689_ _20688_/X VGND VGND VPWR VPWR _20689_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12436__A _12285_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22852__B _22818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13314_/A _13223_/X _13230_/C VGND VGND VPWR VPWR _13231_/C sky130_fd_sc_hd__or3_4
X_25216_ _25219_/CLK _14088_/X HRESETn VGND VGND VPWR VPWR _25216_/Q sky130_fd_sc_hd__dfrtp_4
X_22428_ _22425_/X _22427_/X VGND VGND VPWR VPWR _22428_/Y sky130_fd_sc_hd__nor2_4
XFILLER_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14382__A2 _14380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13161_ _17453_/A VGND VGND VPWR VPWR _13162_/A sky130_fd_sc_hd__inv_2
XANTENNA__15747__A HWDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25147_ _25141_/CLK _25147_/D HRESETn VGND VGND VPWR VPWR _25147_/Q sky130_fd_sc_hd__dfrtp_4
X_22359_ _22355_/X _22358_/X _21767_/X VGND VGND VPWR VPWR _22359_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_108_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14651__A _18010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12112_ _12111_/Y _12107_/X _11842_/X _12107_/X VGND VGND VPWR VPWR _12112_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13092_ _13092_/A _13092_/B VGND VGND VPWR VPWR _13093_/C sky130_fd_sc_hd__nand2_4
X_25078_ _25081_/CLK _14595_/X HRESETn VGND VGND VPWR VPWR _13576_/A sky130_fd_sc_hd__dfrtp_4
X_12043_ _25476_/Q VGND VGND VPWR VPWR _12043_/Y sky130_fd_sc_hd__inv_2
X_16920_ _24247_/Q VGND VGND VPWR VPWR _16920_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13267__A _13457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24029_ _24035_/CLK _24029_/D HRESETn VGND VGND VPWR VPWR _21209_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22601__B1 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24035__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_124_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_124_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16851_ _16850_/Y _16848_/X _16787_/X _16848_/X VGND VGND VPWR VPWR _24404_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15802_ _15809_/A VGND VGND VPWR VPWR _15802_/X sky130_fd_sc_hd__buf_2
X_19570_ _19569_/Y _19567_/X _11943_/X _19567_/X VGND VGND VPWR VPWR _19570_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16782_ _16781_/X VGND VGND VPWR VPWR _16782_/X sky130_fd_sc_hd__buf_2
X_13994_ _13993_/X VGND VGND VPWR VPWR _13995_/B sky130_fd_sc_hd__inv_2
XFILLER_105_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18521_ _18521_/A VGND VGND VPWR VPWR _18541_/A sky130_fd_sc_hd__buf_2
XFILLER_59_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24108__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15733_ _12526_/Y _15732_/X _11778_/X _15732_/X VGND VGND VPWR VPWR _24863_/D sky130_fd_sc_hd__a2bb2o_4
X_12945_ _12945_/A VGND VGND VPWR VPWR _12945_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18452_ _18743_/C VGND VGND VPWR VPWR _18772_/A sky130_fd_sc_hd__buf_2
XFILLER_46_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15664_ _21030_/A VGND VGND VPWR VPWR _15665_/A sky130_fd_sc_hd__buf_2
X_12876_ _12876_/A VGND VGND VPWR VPWR _12876_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17403_ _17403_/A VGND VGND VPWR VPWR _17404_/A sky130_fd_sc_hd__buf_2
X_14615_ _21958_/A VGND VGND VPWR VPWR _14615_/Y sky130_fd_sc_hd__inv_2
X_11827_ _11824_/Y _11816_/X _11825_/X _11826_/X VGND VGND VPWR VPWR _11827_/X sky130_fd_sc_hd__a2bb2o_4
X_18383_ _18383_/A VGND VGND VPWR VPWR _18383_/Y sky130_fd_sc_hd__inv_2
X_15595_ _15595_/A VGND VGND VPWR VPWR _15595_/Y sky130_fd_sc_hd__inv_2
XPHY_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17252_/B _17307_/X _17279_/X _17331_/B VGND VGND VPWR VPWR _17334_/X sky130_fd_sc_hd__a211o_4
XPHY_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11756_/Y _11751_/X _11757_/X _11751_/X VGND VGND VPWR VPWR _11758_/X sky130_fd_sc_hd__a2bb2o_4
X_14546_ _23953_/Q _14546_/B VGND VGND VPWR VPWR _14547_/D sky130_fd_sc_hd__and2_4
XFILLER_81_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_62_0_HCLK clkbuf_8_63_0_HCLK/A VGND VGND VPWR VPWR _24715_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17265_ _17264_/Y _17262_/A VGND VGND VPWR VPWR _17266_/C sky130_fd_sc_hd__or2_4
X_11689_ _25268_/Q VGND VGND VPWR VPWR _11689_/Y sky130_fd_sc_hd__inv_2
X_14477_ _14474_/Y _14476_/X _14411_/X _14476_/X VGND VGND VPWR VPWR _25108_/D sky130_fd_sc_hd__a2bb2o_4
X_19004_ _23879_/Q VGND VGND VPWR VPWR _19004_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24876__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16216_ _16216_/A VGND VGND VPWR VPWR _16216_/Y sky130_fd_sc_hd__inv_2
X_13428_ _13428_/A _13426_/X _13428_/C VGND VGND VPWR VPWR _13428_/X sky130_fd_sc_hd__and3_4
XFILLER_31_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21659__A _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17196_ _17196_/A VGND VGND VPWR VPWR _17196_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17856__B _17846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24805__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13359_ _13455_/A _19717_/A VGND VGND VPWR VPWR _13361_/B sky130_fd_sc_hd__or2_4
X_16147_ HWDATA[8] VGND VGND VPWR VPWR _16147_/X sky130_fd_sc_hd__buf_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16078_ _11739_/A _15646_/A _15927_/X _21053_/A _16077_/X VGND VGND VPWR VPWR _24702_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_116_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15029_ _14966_/A _15027_/Y _25001_/Q _15028_/Y VGND VGND VPWR VPWR _15029_/X sky130_fd_sc_hd__a2bb2o_4
X_19906_ _19906_/A VGND VGND VPWR VPWR _21168_/B sky130_fd_sc_hd__inv_2
XANTENNA__23282__A2_N _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19837_ _19835_/Y _19836_/X _19794_/X _19836_/X VGND VGND VPWR VPWR _23591_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16488__A _24554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19768_ _13426_/B VGND VGND VPWR VPWR _19768_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14833__B1 _25186_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18719_ _18719_/A _18724_/B VGND VGND VPWR VPWR _18721_/B sky130_fd_sc_hd__or2_4
Xclkbuf_5_29_0_HCLK clkbuf_4_14_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19699_ _19699_/A VGND VGND VPWR VPWR _19699_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19772__B1 _19771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21730_ _22923_/A VGND VGND VPWR VPWR _22524_/A sky130_fd_sc_hd__buf_2
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21841__B _22111_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16586__B1 _16228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21661_ _21469_/A _21661_/B _21661_/C VGND VGND VPWR VPWR _21661_/X sky130_fd_sc_hd__or3_4
XFILLER_80_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23400_ _24923_/CLK _23400_/D VGND VGND VPWR VPWR _23400_/Q sky130_fd_sc_hd__dfxtp_4
X_20612_ _15473_/Y _20605_/X _20662_/A _20611_/X VGND VGND VPWR VPWR _20612_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16338__B1 _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24380_ _24391_/CLK _17099_/Y HRESETn VGND VGND VPWR VPWR _17007_/A sky130_fd_sc_hd__dfrtp_4
X_21592_ _21546_/Y _21569_/X _21578_/Y _21592_/D VGND VGND VPWR VPWR _21592_/X sky130_fd_sc_hd__or4_4
XFILLER_32_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23331_ _22795_/A _23322_/Y _23331_/C _23331_/D VGND VGND VPWR VPWR _23331_/X sky130_fd_sc_hd__or4_4
X_20543_ _18871_/X _20542_/Y _20558_/C VGND VGND VPWR VPWR _20543_/X sky130_fd_sc_hd__and3_4
XANTENNA__16889__B2 _16880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12375__A2_N _24837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23084__B1 _22090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23262_ _22820_/X _23262_/B VGND VGND VPWR VPWR _23262_/Y sky130_fd_sc_hd__nor2_4
X_20474_ _14279_/A _20474_/B _24073_/Q VGND VGND VPWR VPWR _20519_/A sky130_fd_sc_hd__and3_4
XANTENNA__19827__B2 _19824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24546__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25001_ _25001_/CLK _15271_/X HRESETn VGND VGND VPWR VPWR _25001_/Q sky130_fd_sc_hd__dfrtp_4
X_22213_ _22193_/X _19246_/Y VGND VGND VPWR VPWR _22214_/C sky130_fd_sc_hd__or2_4
XANTENNA__12375__B2 _24837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21634__A1 _21614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23193_ _23191_/X _23192_/X _22132_/A VGND VGND VPWR VPWR _23193_/X sky130_fd_sc_hd__or3_4
XFILLER_69_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22144_ _22144_/A _22654_/A VGND VGND VPWR VPWR _22144_/X sky130_fd_sc_hd__or2_4
XANTENNA__14190__B _14190_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22075_ _21886_/A _22075_/B VGND VGND VPWR VPWR _22075_/X sky130_fd_sc_hd__or2_4
XFILLER_87_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21026_ _24772_/Q _21026_/B VGND VGND VPWR VPWR _21026_/X sky130_fd_sc_hd__or2_4
XFILLER_102_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18263__B1 _16782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16398__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17530__A1_N _11811_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23008__B _21048_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25334__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22977_ _22975_/X _22976_/X _22485_/X _11776_/A _22775_/X VGND VGND VPWR VPWR _22977_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_43_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12730_ _12731_/A _12731_/B VGND VGND VPWR VPWR _12730_/Y sky130_fd_sc_hd__nand2_4
X_24716_ _24345_/CLK _24716_/D HRESETn VGND VGND VPWR VPWR _16042_/A sky130_fd_sc_hd__dfrtp_4
X_21928_ _21663_/A VGND VGND VPWR VPWR _21929_/A sky130_fd_sc_hd__buf_2
XFILLER_76_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12661_ _12619_/X _12629_/X _12620_/B VGND VGND VPWR VPWR _12662_/C sky130_fd_sc_hd__o21a_4
XFILLER_19_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _15027_/A _21859_/B _21859_/C VGND VGND VPWR VPWR _21859_/X sky130_fd_sc_hd__and3_4
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24647_ _24581_/CLK _24647_/D HRESETn VGND VGND VPWR VPWR _24647_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14646__A _18087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22114__A2 _21548_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18118__A _18221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _16720_/A VGND VGND VPWR VPWR _14400_/X sky130_fd_sc_hd__buf_2
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12592_/A VGND VGND VPWR VPWR _12623_/A sky130_fd_sc_hd__inv_2
X_15380_ _15128_/Y _15379_/X VGND VGND VPWR VPWR _15380_/X sky130_fd_sc_hd__or2_4
XFILLER_19_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24578_ _24596_/CLK _16427_/X HRESETn VGND VGND VPWR VPWR _24578_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22863__A _22186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ _25155_/Q _14330_/X _14327_/A VGND VGND VPWR VPWR _14331_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_7_49_0_HCLK clkbuf_6_24_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_99_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11810__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23529_ _24923_/CLK _23529_/D VGND VGND VPWR VPWR _23529_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _14261_/Y _14259_/X _13837_/X _14259_/X VGND VGND VPWR VPWR _25178_/D sky130_fd_sc_hd__a2bb2o_4
X_17050_ _17050_/A _16981_/Y _17060_/A _17050_/D VGND VGND VPWR VPWR _17051_/B sky130_fd_sc_hd__or4_4
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24287__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13213_ _13227_/A VGND VGND VPWR VPWR _13373_/A sky130_fd_sc_hd__buf_2
X_16001_ _24732_/Q VGND VGND VPWR VPWR _16001_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15477__A _15986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23949__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14193_ _14192_/X VGND VGND VPWR VPWR _14194_/A sky130_fd_sc_hd__buf_2
XANTENNA__22822__B1 _17758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14381__A _14381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24216__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13144_ _24191_/Q VGND VGND VPWR VPWR _13233_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13075_ _12352_/Y _13073_/A VGND VGND VPWR VPWR _13075_/X sky130_fd_sc_hd__or2_4
X_17952_ _17955_/A _19398_/A VGND VGND VPWR VPWR _17952_/X sky130_fd_sc_hd__or2_4
XANTENNA__13866__A1 _20663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12026_ _12013_/X _12018_/X _12026_/C _12026_/D VGND VGND VPWR VPWR _12026_/X sky130_fd_sc_hd__or4_4
X_16903_ _16165_/Y _21048_/A _16165_/Y _21048_/A VGND VGND VPWR VPWR _16904_/D sky130_fd_sc_hd__a2bb2o_4
X_17883_ _16927_/X _17848_/B VGND VGND VPWR VPWR _17883_/Y sky130_fd_sc_hd__nand2_4
XFILLER_120_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19622_ _19622_/A VGND VGND VPWR VPWR _19622_/X sky130_fd_sc_hd__buf_2
X_16834_ _24413_/Q VGND VGND VPWR VPWR _16834_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16101__A _16094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19553_ _11856_/X VGND VGND VPWR VPWR _19553_/X sky130_fd_sc_hd__buf_2
XANTENNA__21942__A _21942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16765_ _16763_/Y _16759_/X _15745_/X _16764_/X VGND VGND VPWR VPWR _24447_/D sky130_fd_sc_hd__a2bb2o_4
X_13977_ _25220_/Q VGND VGND VPWR VPWR _13977_/X sky130_fd_sc_hd__buf_2
XANTENNA__25075__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18504_ _18517_/A _18504_/B _18504_/C VGND VGND VPWR VPWR _18504_/X sky130_fd_sc_hd__and3_4
X_15716_ _15740_/A VGND VGND VPWR VPWR _15763_/A sky130_fd_sc_hd__inv_2
XFILLER_4_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15940__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12928_ _12936_/A _12928_/B _12927_/X VGND VGND VPWR VPWR _25370_/D sky130_fd_sc_hd__and3_4
X_19484_ _19482_/Y _19483_/X _11952_/X _19483_/X VGND VGND VPWR VPWR _23711_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16568__B1 _16398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25004__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16696_ _22560_/A _16695_/X _16340_/X _16695_/X VGND VGND VPWR VPWR _24476_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18435_ _16227_/Y _24160_/Q _16227_/Y _24160_/Q VGND VGND VPWR VPWR _18436_/D sky130_fd_sc_hd__a2bb2o_4
X_15647_ _11865_/X VGND VGND VPWR VPWR _15647_/X sky130_fd_sc_hd__buf_2
XFILLER_62_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12859_ _12859_/A _12858_/Y VGND VGND VPWR VPWR _12861_/B sky130_fd_sc_hd__or2_4
XANTENNA__22105__A2 _22104_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23302__A1 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18028__A _17996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23302__B2 _22833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18366_ _18355_/A _18352_/Y _18365_/X _24187_/Q _18355_/Y VGND VGND VPWR VPWR _18366_/X
+ sky130_fd_sc_hd__a32o_4
X_15578_ _15577_/Y _15575_/X _11767_/X _15575_/X VGND VGND VPWR VPWR _15578_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22656__A3 _22130_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17317_ _17254_/A _17203_/Y _17253_/Y _17320_/B VGND VGND VPWR VPWR _17323_/B sky130_fd_sc_hd__or4_4
X_14529_ _14521_/X _14528_/X _25103_/Q _14517_/A VGND VGND VPWR VPWR _25091_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11801__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18297_ _21491_/A _18296_/X _21491_/A _18296_/X VGND VGND VPWR VPWR _18297_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17248_ _17248_/A VGND VGND VPWR VPWR _22659_/A sky130_fd_sc_hd__inv_2
XANTENNA__16740__B1 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15543__B2 _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_6_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17179_ _22971_/A _17252_/C _24626_/Q _17178_/Y VGND VGND VPWR VPWR _17179_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20190_ _20189_/X VGND VGND VPWR VPWR _20203_/A sky130_fd_sc_hd__inv_2
XANTENNA__18698__A _18705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21836__B _22927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23939__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11868__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19993__B1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22900_ _22770_/X _22899_/X _22479_/X _24722_/Q _22480_/X VGND VGND VPWR VPWR _22900_/X
+ sky130_fd_sc_hd__a32o_4
X_23880_ _23884_/CLK _19003_/X VGND VGND VPWR VPWR _23880_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_110_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21274__D _21273_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22831_ _22520_/A VGND VGND VPWR VPWR _22832_/B sky130_fd_sc_hd__buf_2
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15850__A _15713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21571__B _22835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22762_ _22759_/X _22760_/X _22466_/X _24823_/Q _22761_/X VGND VGND VPWR VPWR _22763_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16559__B1 _16297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21713_ _21331_/X _21713_/B VGND VGND VPWR VPWR _21713_/Y sky130_fd_sc_hd__nor2_4
X_24501_ _23467_/CLK _24501_/D HRESETn VGND VGND VPWR VPWR _13740_/A sky130_fd_sc_hd__dfrtp_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25481_ _25284_/CLK _25481_/D HRESETn VGND VGND VPWR VPWR _25481_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21290__C _21290_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ _22693_/A VGND VGND VPWR VPWR _22693_/Y sky130_fd_sc_hd__inv_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24798__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21644_ _18272_/A _21641_/X _21502_/A _21643_/Y VGND VGND VPWR VPWR _21645_/A sky130_fd_sc_hd__a211o_4
XANTENNA__12045__B1 _25475_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24432_ _25002_/CLK _16798_/X HRESETn VGND VGND VPWR VPWR _24432_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22683__A _23126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24727__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24363_ _24362_/CLK _24363_/D HRESETn VGND VGND VPWR VPWR _17039_/A sky130_fd_sc_hd__dfrtp_4
X_21575_ _16535_/Y _22695_/C VGND VGND VPWR VPWR _21575_/X sky130_fd_sc_hd__and2_4
XFILLER_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15901__A1_N _12769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23314_ _23314_/A _23314_/B VGND VGND VPWR VPWR _23314_/X sky130_fd_sc_hd__and2_4
X_20526_ _20488_/B _20468_/Y _20483_/B _20525_/X VGND VGND VPWR VPWR _20526_/X sky130_fd_sc_hd__a211o_4
XFILLER_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21299__A _23097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24294_ _25433_/CLK _17646_/X HRESETn VGND VGND VPWR VPWR _24294_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16731__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24380__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12348__B2 _24819_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23245_ _22808_/X _23245_/B _23245_/C VGND VGND VPWR VPWR _23245_/X sky130_fd_sc_hd__and3_4
X_20457_ _20496_/C _20452_/X _20420_/B _20457_/D VGND VGND VPWR VPWR _20458_/D sky130_fd_sc_hd__and4_4
XFILLER_4_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22804__B1 _22524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23189__A2_N _23186_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23176_ _23208_/A _23176_/B _23169_/X _23176_/D VGND VGND VPWR VPWR _23176_/X sky130_fd_sc_hd__or4_4
X_20388_ _23384_/Q VGND VGND VPWR VPWR _21969_/A sky130_fd_sc_hd__inv_2
XFILLER_134_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20291__B1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22127_ _21287_/Y _22124_/X _22127_/C VGND VGND VPWR VPWR _22127_/X sky130_fd_sc_hd__and3_4
XANTENNA__18401__A _24172_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22058_ _22053_/X _22057_/X _21767_/X VGND VGND VPWR VPWR _22058_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__11859__B1 _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25515__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13900_ _13899_/X VGND VGND VPWR VPWR _13905_/A sky130_fd_sc_hd__inv_2
X_21009_ _15701_/B VGND VGND VPWR VPWR _21009_/X sky130_fd_sc_hd__buf_2
X_14880_ _14870_/A _14880_/B VGND VGND VPWR VPWR _14880_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__16798__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21791__B1 _17722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21762__A _21618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13831_ _13831_/A VGND VGND VPWR VPWR _13831_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18858__A1_N _16485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22577__B _22727_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12267__A2_N _24765_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16550_ _16550_/A VGND VGND VPWR VPWR _16558_/A sky130_fd_sc_hd__buf_2
XANTENNA__19232__A _16786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13762_ _13762_/A VGND VGND VPWR VPWR _13762_/X sky130_fd_sc_hd__buf_2
Xclkbuf_5_12_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__21543__B1 _14169_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15501_ _11727_/B VGND VGND VPWR VPWR _15501_/Y sky130_fd_sc_hd__inv_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12713_ _12698_/A _12713_/B _12712_/Y VGND VGND VPWR VPWR _25398_/D sky130_fd_sc_hd__and3_4
XFILLER_71_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16481_ _24557_/Q VGND VGND VPWR VPWR _16481_/Y sky130_fd_sc_hd__inv_2
X_13693_ _13693_/A _13693_/B _13693_/C _13693_/D VGND VGND VPWR VPWR _13693_/X sky130_fd_sc_hd__and4_4
XFILLER_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18220_ _18220_/A _18218_/X _18220_/C VGND VGND VPWR VPWR _18224_/B sky130_fd_sc_hd__and3_4
X_15432_ _15446_/A VGND VGND VPWR VPWR _15432_/X sky130_fd_sc_hd__buf_2
X_12644_ _25415_/Q _12644_/B VGND VGND VPWR VPWR _12644_/X sky130_fd_sc_hd__or2_4
XANTENNA__23296__B1 _23172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24468__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18151_ _18215_/A _23879_/Q VGND VGND VPWR VPWR _18152_/C sky130_fd_sc_hd__or2_4
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ _12683_/A _12559_/A _25409_/Q _12526_/Y VGND VGND VPWR VPWR _12575_/X sky130_fd_sc_hd__a2bb2o_4
X_15363_ _15296_/A _15362_/X _15339_/X VGND VGND VPWR VPWR _15363_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_54_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17102_ _17034_/A _17034_/B _17105_/A _17105_/B VGND VGND VPWR VPWR _17108_/B sky130_fd_sc_hd__or4_4
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314_ _14306_/X _14313_/X _13481_/A _14311_/X VGND VGND VPWR VPWR _25163_/D sky130_fd_sc_hd__o22a_4
X_18082_ _18000_/A _18082_/B _18082_/C VGND VGND VPWR VPWR _18086_/B sky130_fd_sc_hd__and3_4
XANTENNA__25088__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15294_ _15080_/Y _15338_/A VGND VGND VPWR VPWR _15307_/C sky130_fd_sc_hd__or2_4
XFILLER_11_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17033_ _16972_/Y _17105_/A _17033_/C _17033_/D VGND VGND VPWR VPWR _17033_/X sky130_fd_sc_hd__or4_4
X_14245_ _13917_/X _14244_/X VGND VGND VPWR VPWR _14245_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_136_0_HCLK clkbuf_7_68_0_HCLK/X VGND VGND VPWR VPWR _23772_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24050__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14176_ _14176_/A VGND VGND VPWR VPWR _25199_/D sky130_fd_sc_hd__inv_2
XANTENNA__21937__A _17717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_199_0_HCLK clkbuf_7_99_0_HCLK/X VGND VGND VPWR VPWR _24909_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_113_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13127_ _20699_/A _13127_/B VGND VGND VPWR VPWR _13128_/B sky130_fd_sc_hd__or2_4
XANTENNA__19407__A _18996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18984_ _23885_/Q VGND VGND VPWR VPWR _18984_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13058_ _13061_/A _13064_/B VGND VGND VPWR VPWR _13062_/B sky130_fd_sc_hd__or2_4
X_17935_ _14648_/X _17933_/X _17934_/X VGND VGND VPWR VPWR _17935_/X sky130_fd_sc_hd__and3_4
XANTENNA__23220__B1 _11753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25256__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12009_ _24088_/Q _11992_/X _12008_/Y VGND VGND VPWR VPWR _12010_/A sky130_fd_sc_hd__o21a_4
XFILLER_61_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12511__B2 _24853_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17866_ _16928_/Y _17850_/D VGND VGND VPWR VPWR _17867_/B sky130_fd_sc_hd__or2_4
XFILLER_93_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16789__B1 _16442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16817_ _14904_/Y _16816_/X HWDATA[21] _16816_/X VGND VGND VPWR VPWR _16817_/X sky130_fd_sc_hd__a2bb2o_4
X_19605_ _19604_/Y _19602_/X _19462_/X _19602_/X VGND VGND VPWR VPWR _23670_/D sky130_fd_sc_hd__a2bb2o_4
X_17797_ _17743_/A _17794_/X VGND VGND VPWR VPWR _17798_/C sky130_fd_sc_hd__or2_4
XFILLER_81_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19536_ _19535_/X VGND VGND VPWR VPWR _19536_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15670__A _15670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16748_ _16747_/Y _16743_/X _16398_/X _16743_/X VGND VGND VPWR VPWR _16748_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21534__B1 _24705_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19467_ _18280_/X VGND VGND VPWR VPWR _20338_/B sky130_fd_sc_hd__buf_2
X_16679_ _16678_/Y _16676_/X _16410_/X _16676_/X VGND VGND VPWR VPWR _16679_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24891__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18418_ _24147_/Q VGND VGND VPWR VPWR _18418_/Y sky130_fd_sc_hd__inv_2
X_19398_ _19398_/A VGND VGND VPWR VPWR _19398_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22629__A3 _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24820__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18349_ _18348_/Y _17478_/X _24188_/Q _17482_/X VGND VGND VPWR VPWR _18363_/A sky130_fd_sc_hd__o22a_4
XFILLER_72_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24138__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21360_ _21547_/A _21360_/B VGND VGND VPWR VPWR _21360_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_7_32_0_HCLK clkbuf_7_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_65_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16713__B1 _16359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22904__A2_N _22901_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20311_ _20298_/Y VGND VGND VPWR VPWR _20311_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_95_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21291_ _21098_/A VGND VGND VPWR VPWR _22705_/A sky130_fd_sc_hd__buf_2
XANTENNA__22950__B _23019_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23030_ _23007_/X _23030_/B _23030_/C _23030_/D VGND VGND VPWR VPWR HRDATA[22] sky130_fd_sc_hd__or4_4
X_20242_ _13341_/B VGND VGND VPWR VPWR _20242_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22262__A1 _21270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20908__A1_N _20882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15845__A _15845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20173_ _20172_/Y _20170_/X _20082_/X _20170_/X VGND VGND VPWR VPWR _20173_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18221__A _18221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_HCLK clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24981_ _24980_/CLK _24981_/D HRESETn VGND VGND VPWR VPWR _24981_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23932_ _25122_/CLK _23932_/D HRESETn VGND VGND VPWR VPWR _20537_/B sky130_fd_sc_hd__dfrtp_4
X_23863_ _25488_/CLK _23863_/D VGND VGND VPWR VPWR _23863_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16676__A _16664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19718__B1 _19599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24979__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22814_ _22808_/X _22814_/B _22814_/C VGND VGND VPWR VPWR _22814_/X sky130_fd_sc_hd__and3_4
XFILLER_72_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23794_ _24396_/CLK _23794_/D VGND VGND VPWR VPWR _23794_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_129_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24908__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25533_ _24692_/CLK _11762_/X HRESETn VGND VGND VPWR VPWR _25533_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22745_ _22745_/A _23035_/A VGND VGND VPWR VPWR _22745_/X sky130_fd_sc_hd__or2_4
XFILLER_26_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23005__C _23005_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25464_ _24383_/CLK _12105_/X HRESETn VGND VGND VPWR VPWR _25464_/Q sky130_fd_sc_hd__dfrtp_4
X_22676_ _15604_/Y _22913_/A VGND VGND VPWR VPWR _22676_/X sky130_fd_sc_hd__and2_4
XANTENNA__24561__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21627_ _21623_/A _20056_/Y VGND VGND VPWR VPWR _21628_/C sky130_fd_sc_hd__or2_4
XFILLER_51_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24415_ _24413_/CLK _16831_/X HRESETn VGND VGND VPWR VPWR _24415_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21828__B2 _22677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25395_ _25397_/CLK _25395_/D HRESETn VGND VGND VPWR VPWR _25395_/Q sky130_fd_sc_hd__dfrtp_4
X_12360_ _12353_/X _12355_/X _12360_/C _12359_/X VGND VGND VPWR VPWR _12381_/B sky130_fd_sc_hd__or4_4
X_21558_ _21556_/X _21558_/B VGND VGND VPWR VPWR _21558_/X sky130_fd_sc_hd__and2_4
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23021__B _23021_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24346_ _24346_/CLK _24346_/D HRESETn VGND VGND VPWR VPWR _24346_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13518__B1 _13472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20509_ _20517_/D _20508_/X VGND VGND VPWR VPWR _24071_/D sky130_fd_sc_hd__or2_4
XFILLER_126_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12291_ _12291_/A _12290_/X VGND VGND VPWR VPWR _12391_/A sky130_fd_sc_hd__or2_4
XFILLER_107_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24277_ _24288_/CLK _24277_/D HRESETn VGND VGND VPWR VPWR _21686_/A sky130_fd_sc_hd__dfrtp_4
X_21489_ _21452_/A _21487_/X _21489_/C VGND VGND VPWR VPWR _21489_/X sky130_fd_sc_hd__and3_4
XANTENNA__12444__A _12286_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14030_ _14030_/A _14030_/B _14001_/X _14040_/D VGND VGND VPWR VPWR _14031_/A sky130_fd_sc_hd__or4_4
XFILLER_88_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22860__B _22626_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_209_0_HCLK clkbuf_7_104_0_HCLK/X VGND VGND VPWR VPWR _24435_/CLK sky130_fd_sc_hd__clkbuf_1
X_23228_ _23119_/X _23226_/X _23121_/X _23227_/X VGND VGND VPWR VPWR _23229_/B sky130_fd_sc_hd__o22a_4
XANTENNA__21757__A _21612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19227__A _19221_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23159_ _16655_/Y _22914_/B VGND VGND VPWR VPWR _23159_/X sky130_fd_sc_hd__and2_4
XFILLER_62_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23202__B1 _22834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15981_ _12181_/Y _15978_/X _15623_/X _15978_/X VGND VGND VPWR VPWR _15981_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17720_ _17719_/Y VGND VGND VPWR VPWR _17720_/X sky130_fd_sc_hd__buf_2
X_14932_ _25004_/Q VGND VGND VPWR VPWR _15063_/A sky130_fd_sc_hd__inv_2
XFILLER_75_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21492__A _21260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17651_ _17651_/A VGND VGND VPWR VPWR _17651_/Y sky130_fd_sc_hd__inv_2
X_14863_ _14824_/X _14862_/Y _14813_/C _14824_/X VGND VGND VPWR VPWR _25032_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16602_ _16599_/Y _16595_/X _16600_/X _16601_/X VGND VGND VPWR VPWR _24511_/D sky130_fd_sc_hd__a2bb2o_4
X_13814_ _14406_/A _15851_/B VGND VGND VPWR VPWR _17413_/A sky130_fd_sc_hd__or2_4
XFILLER_112_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17582_ _17612_/A _17543_/Y _17582_/C _17581_/X VGND VGND VPWR VPWR _17582_/X sky130_fd_sc_hd__or4_4
X_14794_ _13634_/A _13633_/B _14793_/Y _13598_/C _14622_/Y VGND VGND VPWR VPWR _25044_/D
+ sky130_fd_sc_hd__a32o_4
X_19321_ _19320_/Y _19318_/X _19206_/X _19318_/X VGND VGND VPWR VPWR _19321_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24649__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16533_ _24537_/Q VGND VGND VPWR VPWR _16533_/Y sky130_fd_sc_hd__inv_2
X_13745_ _14705_/A VGND VGND VPWR VPWR _13746_/A sky130_fd_sc_hd__buf_2
XFILLER_91_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19252_ _19251_/Y _19249_/X _16876_/X _19249_/X VGND VGND VPWR VPWR _23793_/D sky130_fd_sc_hd__a2bb2o_4
X_16464_ _16463_/Y _16461_/X _16285_/X _16461_/X VGND VGND VPWR VPWR _16464_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15808__A1_N _12368_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13676_ _13676_/A VGND VGND VPWR VPWR _13676_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20836__A _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18203_ _18024_/A _19419_/A VGND VGND VPWR VPWR _18203_/X sky130_fd_sc_hd__or2_4
X_15415_ _15388_/B _15423_/A VGND VGND VPWR VPWR _15415_/X sky130_fd_sc_hd__or2_4
X_12627_ _12657_/A _12625_/X _12626_/X VGND VGND VPWR VPWR _12627_/X sky130_fd_sc_hd__and3_4
X_19183_ _23817_/Q VGND VGND VPWR VPWR _19183_/Y sky130_fd_sc_hd__inv_2
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16395_ _15102_/Y _16389_/X _16393_/X _16394_/X VGND VGND VPWR VPWR _24591_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24231__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18134_ _18023_/X _18132_/X _18134_/C VGND VGND VPWR VPWR _18134_/X sky130_fd_sc_hd__and3_4
X_15346_ _15346_/A _15338_/B _15345_/X VGND VGND VPWR VPWR _24986_/D sky130_fd_sc_hd__and3_4
X_12558_ _12558_/A _12558_/B _12558_/C _12558_/D VGND VGND VPWR VPWR _12558_/X sky130_fd_sc_hd__or4_4
Xclkbuf_6_19_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14553__B HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18065_ _18023_/X _18065_/B _18064_/X VGND VGND VPWR VPWR _18065_/X sky130_fd_sc_hd__and3_4
X_15277_ _15283_/A _15248_/B VGND VGND VPWR VPWR _15278_/B sky130_fd_sc_hd__or2_4
X_12489_ _12209_/Y _12492_/B _12394_/X VGND VGND VPWR VPWR _12489_/Y sky130_fd_sc_hd__a21oi_4
X_17016_ _17016_/A _17013_/X _17014_/X _17016_/D VGND VGND VPWR VPWR _17017_/D sky130_fd_sc_hd__or4_4
X_14228_ _25186_/Q VGND VGND VPWR VPWR _14228_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18448__B1 _16261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14449__A1_N _14169_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25437__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14159_ _14099_/C _14113_/X _14099_/C _14113_/X VGND VGND VPWR VPWR _14159_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18041__A _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18967_ _23892_/Q VGND VGND VPWR VPWR _18967_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25090__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23191__A1_N _12291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17918_ _13541_/A VGND VGND VPWR VPWR _17920_/A sky130_fd_sc_hd__inv_2
X_18898_ _14697_/A VGND VGND VPWR VPWR _19084_/D sky130_fd_sc_hd__buf_2
XFILLER_113_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22498__A _15668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17849_ _17747_/C _17848_/X VGND VGND VPWR VPWR _17850_/D sky130_fd_sc_hd__or2_4
XANTENNA__18620__B1 _16603_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20860_ _20909_/A VGND VGND VPWR VPWR _20860_/X sky130_fd_sc_hd__buf_2
XFILLER_93_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19519_ _22227_/B _19516_/X _11934_/X _19516_/X VGND VGND VPWR VPWR _19519_/X sky130_fd_sc_hd__a2bb2o_4
X_20791_ _20787_/X VGND VGND VPWR VPWR _20791_/Y sky130_fd_sc_hd__inv_2
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24319__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22530_ _22574_/A _22530_/B _22530_/C VGND VGND VPWR VPWR _22530_/X sky130_fd_sc_hd__and3_4
X_22461_ _22786_/A _22460_/X VGND VGND VPWR VPWR _22462_/D sky130_fd_sc_hd__nor2_4
XANTENNA__18216__A _18184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21412_ _21069_/A VGND VGND VPWR VPWR _23034_/A sky130_fd_sc_hd__buf_2
X_24200_ _24305_/CLK _18305_/X HRESETn VGND VGND VPWR VPWR _24200_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22383__D _22383_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25180_ _24955_/CLK _25180_/D HRESETn VGND VGND VPWR VPWR sda_oen_o_S5 sky130_fd_sc_hd__dfstp_4
X_22392_ _21270_/X _22388_/Y _21507_/Y _22391_/X VGND VGND VPWR VPWR _22392_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22961__A _22938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24131_ _24555_/CLK _24131_/D HRESETn VGND VGND VPWR VPWR _24131_/Q sky130_fd_sc_hd__dfrtp_4
X_21343_ _21334_/X _21343_/B _21340_/Y _21343_/D VGND VGND VPWR VPWR _21343_/X sky130_fd_sc_hd__or4_4
XANTENNA__15039__A2_N _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18439__B1 _23232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23954__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24062_ _25397_/CLK _20419_/X HRESETn VGND VGND VPWR VPWR _24062_/Q sky130_fd_sc_hd__dfrtp_4
X_21274_ _21274_/A _21061_/X _21274_/C _21273_/Y VGND VGND VPWR VPWR HRDATA[0] sky130_fd_sc_hd__or4_4
XFILLER_85_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20246__B1 _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23013_ _12252_/Y _22820_/X _23012_/X VGND VGND VPWR VPWR _23013_/Y sky130_fd_sc_hd__o21ai_4
X_20225_ _20223_/Y _20224_/X _19721_/X _20224_/X VGND VGND VPWR VPWR _23447_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15575__A _15563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25107__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_182_0_HCLK clkbuf_7_91_0_HCLK/X VGND VGND VPWR VPWR _25436_/CLK sky130_fd_sc_hd__clkbuf_1
X_20156_ _23473_/Q VGND VGND VPWR VPWR _20156_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24103__D MSI_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_39_0_HCLK clkbuf_8_39_0_HCLK/A VGND VGND VPWR VPWR _25054_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__17790__A _17790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20087_ _20084_/Y _20078_/X _20085_/X _20086_/X VGND VGND VPWR VPWR _23498_/D sky130_fd_sc_hd__a2bb2o_4
X_24964_ _24977_/CLK _24964_/D HRESETn VGND VGND VPWR VPWR _15422_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_135_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24939__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23915_ _24398_/CLK _18905_/X VGND VGND VPWR VPWR _23915_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24895_ _24041_/CLK _24895_/D HRESETn VGND VGND VPWR VPWR _15599_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11860_ _11860_/A VGND VGND VPWR VPWR _11860_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23846_ _23846_/CLK _19101_/X VGND VGND VPWR VPWR _19100_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24742__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11791_ HWDATA[17] VGND VGND VPWR VPWR _11791_/X sky130_fd_sc_hd__buf_2
X_20989_ _14880_/B _20988_/X _20996_/B VGND VGND VPWR VPWR _23988_/D sky130_fd_sc_hd__o21a_4
X_23777_ _23618_/CLK _19298_/X VGND VGND VPWR VPWR _13319_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13530_ _13517_/Y _13529_/Y SCLK_S2 _13529_/A VGND VGND VPWR VPWR _13530_/X sky130_fd_sc_hd__o22a_4
X_25516_ _24285_/CLK _11827_/X HRESETn VGND VGND VPWR VPWR _11824_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_14_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22728_ _22505_/X _22726_/X _21950_/A _22727_/X VGND VGND VPWR VPWR _22728_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17949__B _20209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18390__A2 _17271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13461_ _13461_/A _13461_/B _13460_/X VGND VGND VPWR VPWR _13461_/X sky130_fd_sc_hd__or3_4
X_25447_ _25449_/CLK _25447_/D HRESETn VGND VGND VPWR VPWR _25447_/Q sky130_fd_sc_hd__dfrtp_4
X_22659_ _22659_/A _22534_/X VGND VGND VPWR VPWR _22659_/X sky130_fd_sc_hd__or2_4
X_15200_ _15194_/A _15204_/B _15199_/X _15195_/Y VGND VGND VPWR VPWR _15201_/A sky130_fd_sc_hd__a211o_4
X_12412_ _12412_/A _12407_/B _12411_/X VGND VGND VPWR VPWR _12413_/A sky130_fd_sc_hd__or3_4
X_16180_ _12050_/X _11719_/B _15700_/C _16369_/D VGND VGND VPWR VPWR _16180_/X sky130_fd_sc_hd__or4_4
XANTENNA__12411__B1 _12290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13392_ _13392_/A _13392_/B VGND VGND VPWR VPWR _13392_/X sky130_fd_sc_hd__or2_4
XFILLER_16_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25378_ _25368_/CLK _12897_/X HRESETn VGND VGND VPWR VPWR _12896_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_51_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15131_ _15130_/Y _24581_/Q _15130_/Y _24581_/Q VGND VGND VPWR VPWR _15131_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_51_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12343_ _25339_/Q _12341_/Y _12995_/A _12345_/A VGND VGND VPWR VPWR _12343_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17965__A _14645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24329_ _24330_/CLK _17383_/X HRESETn VGND VGND VPWR VPWR _24329_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_103_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22590__B _22590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12274_ _12390_/B VGND VGND VPWR VPWR _12509_/A sky130_fd_sc_hd__buf_2
X_15062_ _14975_/Y _15278_/A _15283_/A VGND VGND VPWR VPWR _15248_/A sky130_fd_sc_hd__or3_4
XANTENNA__25530__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14013_ _14040_/D _14012_/X VGND VGND VPWR VPWR _14013_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15485__A HTRANS[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19870_ _23579_/Q VGND VGND VPWR VPWR _19870_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12902__A _22660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18821_ _18614_/X _18821_/B VGND VGND VPWR VPWR _18822_/C sky130_fd_sc_hd__or2_4
XFILLER_136_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18752_ _18752_/A VGND VGND VPWR VPWR _18752_/Y sky130_fd_sc_hd__inv_2
X_15964_ HWDATA[17] VGND VGND VPWR VPWR _15964_/X sky130_fd_sc_hd__buf_2
XFILLER_76_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17703_ _17735_/B VGND VGND VPWR VPWR _18319_/B sky130_fd_sc_hd__buf_2
XANTENNA__22934__C1 _22933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14915_ _14915_/A VGND VGND VPWR VPWR _15063_/B sky130_fd_sc_hd__inv_2
XFILLER_23_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18683_ _18683_/A _18619_/Y _18607_/Y _18683_/D VGND VGND VPWR VPWR _18683_/X sky130_fd_sc_hd__or4_4
X_15895_ _15705_/X _15894_/X _11818_/A _24783_/Q _15864_/A VGND VGND VPWR VPWR _24783_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_75_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17634_ _17567_/D _17626_/B VGND VGND VPWR VPWR _17635_/B sky130_fd_sc_hd__or2_4
X_14846_ _25037_/Q _14816_/B _25037_/Q _14816_/B VGND VGND VPWR VPWR _14846_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24483__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17565_ _17565_/A VGND VGND VPWR VPWR _17565_/Y sky130_fd_sc_hd__inv_2
X_14777_ _25046_/Q _25045_/Q _13739_/B _14772_/A VGND VGND VPWR VPWR _14778_/A sky130_fd_sc_hd__a211o_4
XFILLER_91_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11989_ _11989_/A VGND VGND VPWR VPWR _11989_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22162__B1 _14128_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19304_ _13419_/B VGND VGND VPWR VPWR _19304_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24412__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16516_ _16504_/A VGND VGND VPWR VPWR _16516_/X sky130_fd_sc_hd__buf_2
XFILLER_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13728_ _13684_/B _13727_/Y _13721_/X _13714_/A _11669_/A VGND VGND VPWR VPWR _25271_/D
+ sky130_fd_sc_hd__a32o_4
X_17496_ _11763_/Y _17562_/A _11763_/Y _17562_/A VGND VGND VPWR VPWR _17497_/D sky130_fd_sc_hd__a2bb2o_4
X_19235_ _19221_/Y VGND VGND VPWR VPWR _19235_/X sky130_fd_sc_hd__buf_2
X_16447_ _16447_/A VGND VGND VPWR VPWR _16448_/A sky130_fd_sc_hd__inv_2
X_13659_ _13659_/A _13659_/B _24038_/Q _20851_/A VGND VGND VPWR VPWR _13659_/X sky130_fd_sc_hd__or4_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19166_ _19166_/A VGND VGND VPWR VPWR _19166_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16378_ _16378_/A VGND VGND VPWR VPWR _16378_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18117_ _18000_/A _18115_/X _18117_/C VGND VGND VPWR VPWR _18121_/B sky130_fd_sc_hd__and3_4
X_15329_ _15329_/A VGND VGND VPWR VPWR _15329_/Y sky130_fd_sc_hd__inv_2
X_19097_ _23847_/Q VGND VGND VPWR VPWR _19097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14155__B1 _25124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18048_ _18185_/A _18048_/B _18048_/C VGND VGND VPWR VPWR _18059_/B sky130_fd_sc_hd__or3_4
XANTENNA__25271__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25200__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20010_ _21926_/B _20007_/X _19985_/X _20007_/X VGND VGND VPWR VPWR _23529_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_255_0_HCLK clkbuf_8_255_0_HCLK/A VGND VGND VPWR VPWR _25400_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_86_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19999_ _19999_/A VGND VGND VPWR VPWR _22333_/B sky130_fd_sc_hd__inv_2
XFILLER_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21728__B1 _21723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21961_ _21962_/A _19598_/A _14613_/Y _23671_/Q VGND VGND VPWR VPWR _21961_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13643__A _13536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23700_ _23683_/CLK _23700_/D VGND VGND VPWR VPWR _19513_/A sky130_fd_sc_hd__dfxtp_4
X_20912_ _20910_/Y _20906_/X _20911_/X VGND VGND VPWR VPWR _20912_/X sky130_fd_sc_hd__o21a_4
X_21892_ _21887_/X _21892_/B VGND VGND VPWR VPWR _21893_/C sky130_fd_sc_hd__or2_4
X_24680_ _24682_/CLK _16136_/X HRESETn VGND VGND VPWR VPWR _22631_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20951__A1 _25313_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16080__B1 _24701_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _16704_/Y _20836_/X _20824_/X _20842_/Y VGND VGND VPWR VPWR _20843_/X sky130_fd_sc_hd__o22a_4
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23631_ _23388_/CLK _23631_/D VGND VGND VPWR VPWR _19719_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20774_ _20747_/A VGND VGND VPWR VPWR _20774_/X sky130_fd_sc_hd__buf_2
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23562_ _23562_/CLK _23562_/D VGND VGND VPWR VPWR _19915_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25301_ _25301_/CLK _25301_/D HRESETn VGND VGND VPWR VPWR _11990_/A sky130_fd_sc_hd__dfrtp_4
X_22513_ _22513_/A _22513_/B VGND VGND VPWR VPWR _22513_/X sky130_fd_sc_hd__and2_4
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23493_ _23494_/CLK _23493_/D VGND VGND VPWR VPWR _20101_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_10_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22444_ _22444_/A VGND VGND VPWR VPWR _22444_/X sky130_fd_sc_hd__buf_2
X_25232_ _24151_/CLK _25232_/D HRESETn VGND VGND VPWR VPWR _25232_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25359__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22375_ _21887_/X _19908_/Y VGND VGND VPWR VPWR _22375_/X sky130_fd_sc_hd__or2_4
X_25163_ _25309_/CLK _25163_/D HRESETn VGND VGND VPWR VPWR _25163_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21326_ _22798_/A VGND VGND VPWR VPWR _21326_/X sky130_fd_sc_hd__buf_2
XFILLER_124_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24114_ _24120_/CLK _18820_/X HRESETn VGND VGND VPWR VPWR _24114_/Q sky130_fd_sc_hd__dfrtp_4
X_25094_ _25137_/CLK _14523_/X HRESETn VGND VGND VPWR VPWR _25094_/Q sky130_fd_sc_hd__dfrtp_4
X_21257_ _21247_/A _21255_/X _21257_/C VGND VGND VPWR VPWR _21257_/X sky130_fd_sc_hd__and3_4
X_24045_ _24413_/CLK _20891_/X HRESETn VGND VGND VPWR VPWR _20889_/A sky130_fd_sc_hd__dfrtp_4
X_20208_ _21231_/B _20203_/X _20123_/X _20203_/A VGND VGND VPWR VPWR _20208_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18832__B1 _16483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21188_ _21186_/A VGND VGND VPWR VPWR _21191_/A sky130_fd_sc_hd__buf_2
XFILLER_81_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13535__A1_N SSn_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24994__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20139_ _20139_/A VGND VGND VPWR VPWR _21629_/B sky130_fd_sc_hd__inv_2
XANTENNA__21982__A3 _21951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24923__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12961_ _12774_/Y _12964_/B _12866_/X VGND VGND VPWR VPWR _12961_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16462__A1_N _16457_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24947_ _24950_/CLK _15459_/X HRESETn VGND VGND VPWR VPWR _13927_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14700_ _21388_/A VGND VGND VPWR VPWR _21614_/A sky130_fd_sc_hd__buf_2
X_11912_ _11878_/B _11902_/B _11916_/B VGND VGND VPWR VPWR _11912_/Y sky130_fd_sc_hd__o21ai_4
X_15680_ _15680_/A VGND VGND VPWR VPWR _15687_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_5_15_0_HCLK_A clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12892_ _12881_/A _12890_/X _12891_/X VGND VGND VPWR VPWR _25380_/D sky130_fd_sc_hd__and3_4
XFILLER_2_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24878_ _24026_/CLK _24878_/D HRESETn VGND VGND VPWR VPWR _20812_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14631_ _14623_/X _14630_/Y _14613_/A _14622_/Y VGND VGND VPWR VPWR _14631_/X sky130_fd_sc_hd__a2bb2o_4
X_11843_ _11840_/Y _11836_/X _11842_/X _11836_/X VGND VGND VPWR VPWR _11843_/X sky130_fd_sc_hd__a2bb2o_4
X_23829_ _25044_/CLK _19150_/X VGND VGND VPWR VPWR _23829_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12176__A1_N _14329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17350_ _17350_/A _17350_/B _17350_/C _17349_/X VGND VGND VPWR VPWR _17353_/B sky130_fd_sc_hd__or4_4
XFILLER_54_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16477__A1_N _16476_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14562_ _13573_/Y _14561_/X VGND VGND VPWR VPWR _14563_/B sky130_fd_sc_hd__or2_4
XFILLER_14_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11774_ HWDATA[22] VGND VGND VPWR VPWR _11774_/X sky130_fd_sc_hd__buf_2
X_16301_ _16299_/Y _16296_/X _16300_/X _16296_/X VGND VGND VPWR VPWR _24624_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13513_ _13511_/Y _13507_/X _11858_/X _13512_/X VGND VGND VPWR VPWR _13513_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17281_ _17280_/X VGND VGND VPWR VPWR _24356_/D sky130_fd_sc_hd__inv_2
X_14493_ _14492_/Y _14488_/X _14400_/X _14481_/A VGND VGND VPWR VPWR _14493_/X sky130_fd_sc_hd__a2bb2o_4
X_19020_ _19020_/A VGND VGND VPWR VPWR _19020_/Y sky130_fd_sc_hd__inv_2
X_16232_ _16225_/A VGND VGND VPWR VPWR _16232_/X sky130_fd_sc_hd__buf_2
XANTENNA__14385__B1 _13835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13444_ _13312_/A _23501_/Q VGND VGND VPWR VPWR _13445_/C sky130_fd_sc_hd__or2_4
XFILLER_70_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16163_ _21426_/A VGND VGND VPWR VPWR _16163_/Y sky130_fd_sc_hd__inv_2
X_13375_ _13173_/X _13371_/X _13374_/X VGND VGND VPWR VPWR _13375_/X sky130_fd_sc_hd__or3_4
XANTENNA__25029__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15114_ _15114_/A VGND VGND VPWR VPWR _15388_/B sky130_fd_sc_hd__inv_2
X_12326_ _12326_/A _12319_/X _12326_/C _12325_/X VGND VGND VPWR VPWR _12340_/C sky130_fd_sc_hd__or4_4
X_16094_ _16094_/A VGND VGND VPWR VPWR _16094_/X sky130_fd_sc_hd__buf_2
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15885__B1 _11791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21010__A _21009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15045_ _15210_/B _24447_/Q _15210_/B _24447_/Q VGND VGND VPWR VPWR _15047_/C sky130_fd_sc_hd__a2bb2o_4
X_19922_ _19922_/A VGND VGND VPWR VPWR _21618_/B sky130_fd_sc_hd__inv_2
X_12257_ _12257_/A VGND VGND VPWR VPWR _12257_/Y sky130_fd_sc_hd__inv_2
X_12188_ _12188_/A VGND VGND VPWR VPWR _12440_/C sky130_fd_sc_hd__buf_2
X_19853_ _19851_/Y _19847_/X _19783_/X _19852_/X VGND VGND VPWR VPWR _19853_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15637__B1 _14470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11910__A2 _11700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18804_ _18623_/Y _18803_/X _18707_/X VGND VGND VPWR VPWR _18804_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_22_0_HCLK clkbuf_8_22_0_HCLK/A VGND VGND VPWR VPWR _24102_/CLK sky130_fd_sc_hd__clkbuf_1
X_16996_ _16044_/Y _24372_/Q _16044_/Y _24372_/Q VGND VGND VPWR VPWR _16996_/X sky130_fd_sc_hd__a2bb2o_4
X_19784_ _19793_/A VGND VGND VPWR VPWR _19784_/X sky130_fd_sc_hd__buf_2
XANTENNA__24664__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_85_0_HCLK clkbuf_7_42_0_HCLK/X VGND VGND VPWR VPWR _24957_/CLK sky130_fd_sc_hd__clkbuf_1
X_15947_ _15930_/X _15935_/X HWDATA[26] _24761_/Q _15933_/X VGND VGND VPWR VPWR _15947_/X
+ sky130_fd_sc_hd__a32o_4
X_18735_ _18734_/X VGND VGND VPWR VPWR _24137_/D sky130_fd_sc_hd__inv_2
XFILLER_97_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18666_ _18661_/X _18666_/B _18666_/C _18665_/X VGND VGND VPWR VPWR _18666_/X sky130_fd_sc_hd__or4_4
XFILLER_37_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15878_ _12824_/Y _15872_/X _11774_/X _15872_/X VGND VGND VPWR VPWR _15878_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16062__B1 _16061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20933__B2 _20913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14829_ _14831_/A _14827_/X _14226_/Y _14828_/X VGND VGND VPWR VPWR _14829_/X sky130_fd_sc_hd__o22a_4
X_17617_ _17617_/A _17617_/B _17617_/C VGND VGND VPWR VPWR _17617_/X sky130_fd_sc_hd__and3_4
X_18597_ _18677_/A VGND VGND VPWR VPWR _18789_/A sky130_fd_sc_hd__buf_2
XFILLER_63_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22495__B _22493_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17548_ _11753_/A _17559_/A _11844_/Y _17576_/A VGND VGND VPWR VPWR _17550_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22686__A1 _22786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22686__B2 _22685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17479_ _21504_/A _17474_/X _17478_/X VGND VGND VPWR VPWR _24311_/D sky130_fd_sc_hd__a21oi_4
X_19218_ _13182_/B VGND VGND VPWR VPWR _19218_/Y sky130_fd_sc_hd__inv_2
X_20490_ _20490_/A _20489_/Y VGND VGND VPWR VPWR _20490_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__25452__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19149_ _17442_/X VGND VGND VPWR VPWR _19149_/X sky130_fd_sc_hd__buf_2
XANTENNA__22989__A2 _22988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22160_ _22159_/X VGND VGND VPWR VPWR _22160_/Y sky130_fd_sc_hd__inv_2
X_21111_ _21018_/A VGND VGND VPWR VPWR _21111_/X sky130_fd_sc_hd__buf_2
XANTENNA__15876__B1 _11767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22091_ _24539_/Q _21026_/B _21326_/X VGND VGND VPWR VPWR _22091_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12542__A _12542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21042_ _22549_/A _21017_/X _21042_/C VGND VGND VPWR VPWR _21274_/A sky130_fd_sc_hd__and3_4
XANTENNA__21855__A _16723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15891__A3 _11803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22610__A1 _24413_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15639__A1_N _15638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15628__B1 _15627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15853__A _15852_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18290__A1 _24198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24801_ _25385_/CLK _15870_/X HRESETn VGND VGND VPWR VPWR _24801_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14469__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22993_ _16485_/A _22879_/X _22798_/X VGND VGND VPWR VPWR _22993_/X sky130_fd_sc_hd__o21a_4
XFILLER_27_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24334__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24732_ _24355_/CLK _16004_/X HRESETn VGND VGND VPWR VPWR _24732_/Q sky130_fd_sc_hd__dfrtp_4
X_21944_ _21944_/A _19569_/Y VGND VGND VPWR VPWR _21944_/X sky130_fd_sc_hd__or2_4
XANTENNA__16053__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20924__B2 _20913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24663_ _24162_/CLK _24663_/D HRESETn VGND VGND VPWR VPWR _23242_/A sky130_fd_sc_hd__dfrtp_4
X_21875_ _21875_/A _21874_/X VGND VGND VPWR VPWR _21875_/X sky130_fd_sc_hd__and2_4
XFILLER_131_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15800__B1 _11749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23623_/CLK _23614_/D VGND VGND VPWR VPWR _13426_/B sky130_fd_sc_hd__dfxtp_4
X_20826_ _21582_/A _20815_/X _20824_/X _20825_/X VGND VGND VPWR VPWR _20827_/A sky130_fd_sc_hd__o22a_4
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24594_ _24596_/CLK _24594_/D HRESETn VGND VGND VPWR VPWR _15090_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23545_ _23545_/CLK _23545_/D VGND VGND VPWR VPWR _23545_/Q sky130_fd_sc_hd__dfxtp_4
X_20757_ _13119_/B VGND VGND VPWR VPWR _20757_/Y sky130_fd_sc_hd__inv_2
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20688_ _21584_/A _20677_/X _20686_/X _20687_/X VGND VGND VPWR VPWR _20688_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23476_ _23516_/CLK _23476_/D VGND VGND VPWR VPWR _23476_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_137_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25193__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25215_ _25219_/CLK _25215_/D HRESETn VGND VGND VPWR VPWR _13985_/B sky130_fd_sc_hd__dfrtp_4
X_22427_ _16146_/Y _22426_/X _22422_/X _11828_/Y _22265_/X VGND VGND VPWR VPWR _22427_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_13_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13160_ _13188_/A _13158_/X _13159_/X VGND VGND VPWR VPWR _13160_/X sky130_fd_sc_hd__and3_4
XFILLER_136_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25146_ _25141_/CLK _25146_/D HRESETn VGND VGND VPWR VPWR _25146_/Q sky130_fd_sc_hd__dfrtp_4
X_22358_ _21885_/X _22356_/X _22357_/X VGND VGND VPWR VPWR _22358_/X sky130_fd_sc_hd__and3_4
XFILLER_123_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12111_ _25461_/Q VGND VGND VPWR VPWR _12111_/Y sky130_fd_sc_hd__inv_2
X_13091_ _13076_/A _13087_/X _13090_/Y VGND VGND VPWR VPWR _13091_/X sky130_fd_sc_hd__and3_4
X_21309_ _16723_/A VGND VGND VPWR VPWR _23170_/A sky130_fd_sc_hd__buf_2
X_22289_ _13658_/A VGND VGND VPWR VPWR _22289_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12452__A _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25077_ _25290_/CLK _25077_/D HRESETn VGND VGND VPWR VPWR _14559_/A sky130_fd_sc_hd__dfrtp_4
X_12042_ _12040_/Y _12041_/X _25476_/Q _12041_/X VGND VGND VPWR VPWR _25477_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24028_ _24909_/CLK _24028_/D HRESETn VGND VGND VPWR VPWR _24028_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16859__A _16880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20612__B1 _20662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16850_ _16850_/A VGND VGND VPWR VPWR _16850_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19235__A _19221_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15801_ _12364_/Y _15799_/X _11754_/X _15799_/X VGND VGND VPWR VPWR _24835_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16292__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16781_ HWDATA[4] VGND VGND VPWR VPWR _16781_/X sky130_fd_sc_hd__buf_2
X_13993_ _14012_/A _14003_/C _14023_/A _13992_/X VGND VGND VPWR VPWR _13993_/X sky130_fd_sc_hd__or4_4
XANTENNA__24075__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18520_ _18520_/A VGND VGND VPWR VPWR _18520_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15732_ _15721_/A VGND VGND VPWR VPWR _15732_/X sky130_fd_sc_hd__buf_2
XFILLER_19_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12944_ _12955_/A _12944_/B _12944_/C _12944_/D VGND VGND VPWR VPWR _12945_/A sky130_fd_sc_hd__or4_4
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19230__B1 _19206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24004__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18451_ _18451_/A _18451_/B VGND VGND VPWR VPWR _18743_/C sky130_fd_sc_hd__or2_4
X_15663_ _15670_/A VGND VGND VPWR VPWR _21030_/A sky130_fd_sc_hd__inv_2
X_12875_ _12840_/Y _12863_/X _12874_/X _12871_/B VGND VGND VPWR VPWR _12876_/A sky130_fd_sc_hd__a211o_4
X_17402_ _23982_/Q _17402_/B VGND VGND VPWR VPWR _17403_/A sky130_fd_sc_hd__or2_4
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14614_ _14613_/Y _13638_/X _14613_/A _13637_/A VGND VGND VPWR VPWR _14614_/X sky130_fd_sc_hd__o22a_4
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11826_ _11794_/X VGND VGND VPWR VPWR _11826_/X sky130_fd_sc_hd__buf_2
X_18382_ _18381_/Y _18377_/X _18383_/A _18377_/X VGND VGND VPWR VPWR _24181_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15594_ _15592_/Y _15588_/X _11788_/X _15593_/X VGND VGND VPWR VPWR _15594_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17333_ _17306_/X _17331_/X _17333_/C VGND VGND VPWR VPWR _24343_/D sky130_fd_sc_hd__and3_4
XANTENNA__19533__B2 _19528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14041_/Y _14049_/X _14545_/C _14054_/Y VGND VGND VPWR VPWR _14546_/B sky130_fd_sc_hd__or4_4
XFILLER_109_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ HWDATA[27] VGND VGND VPWR VPWR _11757_/X sky130_fd_sc_hd__buf_2
XPHY_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17544__B1 _11780_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11752__A2_N _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17264_ _24359_/Q VGND VGND VPWR VPWR _17264_/Y sky130_fd_sc_hd__inv_2
X_14476_ _14481_/A VGND VGND VPWR VPWR _14476_/X sky130_fd_sc_hd__buf_2
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11688_ _11678_/X _11688_/B _11684_/X _11688_/D VGND VGND VPWR VPWR _11688_/X sky130_fd_sc_hd__or4_4
X_19003_ _19002_/Y _18998_/X _18977_/X _18998_/X VGND VGND VPWR VPWR _19003_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16215_ _16214_/Y _16212_/X _15957_/X _16212_/X VGND VGND VPWR VPWR _16215_/X sky130_fd_sc_hd__a2bb2o_4
X_13427_ _13320_/A _19817_/A VGND VGND VPWR VPWR _13428_/C sky130_fd_sc_hd__or2_4
X_17195_ _23247_/A _23246_/A _16287_/Y _17194_/Y VGND VGND VPWR VPWR _17201_/B sky130_fd_sc_hd__o22a_4
X_16146_ _24676_/Q VGND VGND VPWR VPWR _16146_/Y sky130_fd_sc_hd__inv_2
X_13358_ _13390_/A _13358_/B _13357_/X VGND VGND VPWR VPWR _13366_/B sky130_fd_sc_hd__or3_4
X_12309_ _24834_/Q VGND VGND VPWR VPWR _12309_/Y sky130_fd_sc_hd__inv_2
X_16077_ _16079_/A _15843_/A VGND VGND VPWR VPWR _16077_/X sky130_fd_sc_hd__or2_4
X_13289_ _13453_/A _13286_/X _13288_/X VGND VGND VPWR VPWR _13293_/B sky130_fd_sc_hd__and3_4
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24845__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15028_ _24439_/Q VGND VGND VPWR VPWR _15028_/Y sky130_fd_sc_hd__inv_2
X_19905_ _19904_/Y _19902_/X _19632_/X _19902_/X VGND VGND VPWR VPWR _19905_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14530__B1 _21119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16769__A _24444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19836_ _19836_/A VGND VGND VPWR VPWR _19836_/X sky130_fd_sc_hd__buf_2
XFILLER_84_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16283__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19767_ _19765_/Y _19766_/X _19721_/X _19766_/X VGND VGND VPWR VPWR _19767_/X sky130_fd_sc_hd__a2bb2o_4
X_16979_ _24710_/Q _24367_/Q _16056_/Y _17038_/C VGND VGND VPWR VPWR _16980_/D sky130_fd_sc_hd__o22a_4
X_18718_ _18717_/X VGND VGND VPWR VPWR _18724_/B sky130_fd_sc_hd__inv_2
XFILLER_37_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19698_ _19696_/Y _19697_/X _19553_/X _19697_/X VGND VGND VPWR VPWR _23639_/D sky130_fd_sc_hd__a2bb2o_4
X_18649_ _16579_/Y _24130_/Q _24523_/Q _18749_/A VGND VGND VPWR VPWR _18652_/C sky130_fd_sc_hd__a2bb2o_4
X_21660_ _21656_/X _21659_/X _18299_/X VGND VGND VPWR VPWR _21661_/C sky130_fd_sc_hd__o21a_4
XFILLER_51_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20611_ _17388_/X _20609_/Y _20611_/C VGND VGND VPWR VPWR _20611_/X sky130_fd_sc_hd__and3_4
X_21591_ _21103_/X _21586_/Y _21587_/X _21590_/X VGND VGND VPWR VPWR _21592_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16338__B2 _16337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17535__B1 _11776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20542_ _23933_/Q _20539_/A VGND VGND VPWR VPWR _20542_/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23330_ _23207_/A _23327_/X _23330_/C VGND VGND VPWR VPWR _23331_/D sky130_fd_sc_hd__and3_4
XFILLER_20_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23130__A _22798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20473_ _20472_/X VGND VGND VPWR VPWR _20473_/X sky130_fd_sc_hd__buf_2
XANTENNA__15848__A _15674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23261_ _12217_/Y _22426_/X _22712_/X _12328_/Y _22840_/X VGND VGND VPWR VPWR _23262_/B
+ sky130_fd_sc_hd__o32a_4
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14752__A _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18224__A _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25000_ _25001_/CLK _15274_/X HRESETn VGND VGND VPWR VPWR _25000_/Q sky130_fd_sc_hd__dfrtp_4
X_22212_ _21595_/A _22212_/B VGND VGND VPWR VPWR _22212_/X sky130_fd_sc_hd__or2_4
XFILLER_119_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23192_ _17178_/Y _22475_/X _12747_/A _22435_/X VGND VGND VPWR VPWR _23192_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22143_ _22963_/A _22142_/X VGND VGND VPWR VPWR _22143_/X sky130_fd_sc_hd__and2_4
XFILLER_82_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24586__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22074_ _22069_/X _22073_/X _14677_/X VGND VGND VPWR VPWR _22074_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_86_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24515__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21025_ _21025_/A VGND VGND VPWR VPWR _21040_/A sky130_fd_sc_hd__buf_2
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19055__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19460__B1 _19370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16274__B1 _24632_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_HCLK_A clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13815__B _17413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13088__B1 _13031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11830__A1_N _11828_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22976_ _22976_/A _22864_/X VGND VGND VPWR VPWR _22976_/X sky130_fd_sc_hd__or2_4
XFILLER_56_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24715_ _24715_/CLK _16045_/X HRESETn VGND VGND VPWR VPWR _16044_/A sky130_fd_sc_hd__dfrtp_4
X_21927_ _21917_/X _21923_/X _21926_/X VGND VGND VPWR VPWR _21927_/X sky130_fd_sc_hd__and3_4
XFILLER_55_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12660_ _12657_/A _12656_/B _12660_/C VGND VGND VPWR VPWR _12660_/X sky130_fd_sc_hd__and3_4
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24646_ _24581_/CLK _16239_/X HRESETn VGND VGND VPWR VPWR _22619_/A sky130_fd_sc_hd__dfrtp_4
X_21858_ _21323_/A VGND VGND VPWR VPWR _21858_/X sky130_fd_sc_hd__buf_2
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25374__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18443__A1_N _23004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _20807_/Y _20808_/Y _13137_/X VGND VGND VPWR VPWR _20809_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12596_/A _24845_/Q _25389_/Q _12562_/Y VGND VGND VPWR VPWR _12598_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17526__B1 _11840_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24577_ _24596_/CLK _24577_/D HRESETn VGND VGND VPWR VPWR _24577_/Q sky130_fd_sc_hd__dfrtp_4
X_21789_ _21459_/A _21789_/B VGND VGND VPWR VPWR _21789_/X sky130_fd_sc_hd__or2_4
XANTENNA__25303__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _14330_/A VGND VGND VPWR VPWR _14330_/X sky130_fd_sc_hd__buf_2
XFILLER_11_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23528_ _24923_/CLK _20012_/X VGND VGND VPWR VPWR _23528_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20664__A _20664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ _14261_/A VGND VGND VPWR VPWR _14261_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15758__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23459_ _23434_/CLK _20194_/X VGND VGND VPWR VPWR _23459_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16000_ _15999_/Y _15997_/X _11746_/X _15997_/X VGND VGND VPWR VPWR _24733_/D sky130_fd_sc_hd__a2bb2o_4
X_13212_ _13212_/A VGND VGND VPWR VPWR _13227_/A sky130_fd_sc_hd__buf_2
X_14192_ _14192_/A VGND VGND VPWR VPWR _14192_/X sky130_fd_sc_hd__buf_2
XFILLER_136_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13143_ _13177_/A VGND VGND VPWR VPWR _13143_/X sky130_fd_sc_hd__buf_2
XANTENNA__17973__A _17996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25129_ _25113_/CLK _14422_/X HRESETn VGND VGND VPWR VPWR _25129_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__12182__A _25447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13074_ _25335_/Q _13073_/Y VGND VGND VPWR VPWR _13076_/B sky130_fd_sc_hd__or2_4
X_17951_ _17947_/X _17950_/X _18017_/A VGND VGND VPWR VPWR _17951_/X sky130_fd_sc_hd__o21a_4
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24256__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12025_ _12023_/Y _12024_/X _12023_/Y _12024_/X VGND VGND VPWR VPWR _12026_/D sky130_fd_sc_hd__a2bb2o_4
X_16902_ _22976_/A _16900_/Y _23187_/A _17786_/A VGND VGND VPWR VPWR _16904_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17882_ _17874_/A _17878_/X _17882_/C VGND VGND VPWR VPWR _17882_/X sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_5_30_0_HCLK_A clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19621_ _19621_/A VGND VGND VPWR VPWR _19621_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16833_ _16832_/Y _16830_/X _15747_/X _16830_/X VGND VGND VPWR VPWR _16833_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22338__B1 _18298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16764_ _16773_/A VGND VGND VPWR VPWR _16764_/X sky130_fd_sc_hd__buf_2
X_19552_ _19538_/X VGND VGND VPWR VPWR _19552_/X sky130_fd_sc_hd__buf_2
X_13976_ _14036_/A VGND VGND VPWR VPWR _13976_/X sky130_fd_sc_hd__buf_2
XFILLER_19_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12826__B1 _12849_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15715_ _15548_/X _15713_/X _15714_/X _24872_/Q _15711_/X VGND VGND VPWR VPWR _24872_/D
+ sky130_fd_sc_hd__a32o_4
X_18503_ _18503_/A _18503_/B VGND VGND VPWR VPWR _18504_/C sky130_fd_sc_hd__or2_4
XFILLER_74_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12927_ _12927_/A _12927_/B VGND VGND VPWR VPWR _12927_/X sky130_fd_sc_hd__or2_4
XFILLER_98_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16695_ _16645_/A VGND VGND VPWR VPWR _16695_/X sky130_fd_sc_hd__buf_2
X_19483_ _19470_/Y VGND VGND VPWR VPWR _19483_/X sky130_fd_sc_hd__buf_2
XFILLER_111_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_159_0_HCLK clkbuf_7_79_0_HCLK/X VGND VGND VPWR VPWR _24689_/CLK sky130_fd_sc_hd__clkbuf_1
X_15646_ _15646_/A VGND VGND VPWR VPWR _15646_/X sky130_fd_sc_hd__buf_2
X_18434_ _16221_/Y _24162_/Q _22992_/A _18400_/Y VGND VGND VPWR VPWR _18434_/X sky130_fd_sc_hd__a2bb2o_4
X_12858_ _12858_/A VGND VGND VPWR VPWR _12858_/Y sky130_fd_sc_hd__inv_2
X_11809_ _11809_/A VGND VGND VPWR VPWR _11809_/X sky130_fd_sc_hd__buf_2
X_18365_ _18365_/A _18365_/B VGND VGND VPWR VPWR _18365_/X sky130_fd_sc_hd__or2_4
X_15577_ _15577_/A VGND VGND VPWR VPWR _15577_/Y sky130_fd_sc_hd__inv_2
X_12789_ _25357_/Q _24774_/Q _12845_/B _12788_/Y VGND VGND VPWR VPWR _12789_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25044__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17315_/X VGND VGND VPWR VPWR _24348_/D sky130_fd_sc_hd__inv_2
X_14528_ _21542_/A _14510_/X _21334_/A _14505_/X VGND VGND VPWR VPWR _14528_/X sky130_fd_sc_hd__o22a_4
X_18296_ _18300_/A _18295_/Y VGND VGND VPWR VPWR _18296_/X sky130_fd_sc_hd__or2_4
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17247_ _17188_/Y _17169_/A _17243_/X _17247_/D VGND VGND VPWR VPWR _17247_/X sky130_fd_sc_hd__or4_4
X_14459_ _14453_/Y VGND VGND VPWR VPWR _14459_/X sky130_fd_sc_hd__buf_2
XFILLER_128_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17178_ _24355_/Q VGND VGND VPWR VPWR _17178_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22813__A1 _24519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16129_ _16128_/Y _16126_/X _11800_/X _16126_/X VGND VGND VPWR VPWR _16129_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17883__A _16927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19819_ _13459_/B VGND VGND VPWR VPWR _19819_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13635__B _13598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23979__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22830_ _22830_/A VGND VGND VPWR VPWR _22830_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21852__B _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12817__B1 _12843_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_55_0_HCLK clkbuf_7_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16008__B1 _15944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23125__A _22795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22761_ _23097_/A VGND VGND VPWR VPWR _22761_/X sky130_fd_sc_hd__buf_2
XFILLER_112_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13490__B1 _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12293__B2 _24818_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24500_ _23498_/CLK _24500_/D HRESETn VGND VGND VPWR VPWR _13741_/C sky130_fd_sc_hd__dfrtp_4
X_21712_ _21712_/A _21709_/Y _21710_/X _21712_/D VGND VGND VPWR VPWR _21713_/B sky130_fd_sc_hd__and4_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25480_ _25284_/CLK _12035_/X HRESETn VGND VGND VPWR VPWR _12033_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_13_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22692_ _22511_/B _22690_/X _22783_/A _22691_/X VGND VGND VPWR VPWR _22693_/A sky130_fd_sc_hd__o22a_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12045__A1 _24093_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24431_ _24431_/CLK _16800_/X HRESETn VGND VGND VPWR VPWR _16799_/A sky130_fd_sc_hd__dfrtp_4
X_21643_ _21643_/A _21816_/B VGND VGND VPWR VPWR _21643_/Y sky130_fd_sc_hd__nor2_4
XFILLER_40_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22501__B1 _12092_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24362_ _24362_/CLK _17160_/X HRESETn VGND VGND VPWR VPWR _16985_/A sky130_fd_sc_hd__dfrtp_4
X_21574_ _15852_/Y VGND VGND VPWR VPWR _22695_/C sky130_fd_sc_hd__buf_2
XFILLER_36_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23313_ _23281_/A _23313_/B _23313_/C _23312_/X VGND VGND VPWR VPWR _23313_/X sky130_fd_sc_hd__or4_4
X_20525_ _20525_/A _20519_/X VGND VGND VPWR VPWR _20525_/X sky130_fd_sc_hd__and2_4
XFILLER_138_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24293_ _25433_/CLK _17649_/X HRESETn VGND VGND VPWR VPWR _17565_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_101_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24767__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20456_ _20445_/B _20423_/X VGND VGND VPWR VPWR _20457_/D sky130_fd_sc_hd__and2_4
XFILLER_10_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23244_ _24531_/Q _22393_/X _15668_/A _23243_/X VGND VGND VPWR VPWR _23245_/C sky130_fd_sc_hd__a211o_4
XFILLER_119_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20387_ _20385_/Y _20386_/Y _19758_/X _20386_/Y VGND VGND VPWR VPWR _23385_/D sky130_fd_sc_hd__a2bb2o_4
X_23175_ _23207_/A _23175_/B _23174_/X VGND VGND VPWR VPWR _23176_/D sky130_fd_sc_hd__and3_4
XFILLER_137_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23945__D scl_i_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22126_ _22125_/X VGND VGND VPWR VPWR _22127_/C sky130_fd_sc_hd__buf_2
XANTENNA__15837__A3 _15836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22057_ _21885_/X _22054_/X _22056_/X VGND VGND VPWR VPWR _22057_/X sky130_fd_sc_hd__and3_4
XFILLER_134_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23019__B _23019_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21008_ _25286_/Q _21008_/B VGND VGND VPWR VPWR _21008_/X sky130_fd_sc_hd__and2_4
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13830_ _13580_/Y _13829_/X _11822_/X _13829_/X VGND VGND VPWR VPWR _13830_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23035__A _23035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13761_ _13754_/A VGND VGND VPWR VPWR _13762_/A sky130_fd_sc_hd__buf_2
X_22959_ _22958_/X VGND VGND VPWR VPWR _22959_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15500_ _15498_/Y _15499_/X HADDR[19] _15499_/X VGND VGND VPWR VPWR _15500_/X sky130_fd_sc_hd__a2bb2o_4
X_12712_ _12712_/A _12712_/B VGND VGND VPWR VPWR _12712_/Y sky130_fd_sc_hd__nand2_4
X_16480_ _16478_/Y _16474_/X _16393_/X _16479_/X VGND VGND VPWR VPWR _16480_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13692_ _13698_/B VGND VGND VPWR VPWR _13693_/B sky130_fd_sc_hd__inv_2
XFILLER_31_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15431_ _15430_/X VGND VGND VPWR VPWR _15446_/A sky130_fd_sc_hd__buf_2
X_12643_ _12645_/B VGND VGND VPWR VPWR _12644_/B sky130_fd_sc_hd__inv_2
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24629_ _24612_/CLK _24629_/D HRESETn VGND VGND VPWR VPWR _24629_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18150_ _18150_/A _18150_/B VGND VGND VPWR VPWR _18150_/X sky130_fd_sc_hd__or2_4
XFILLER_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15362_ _15367_/A _15369_/A _15365_/A _15365_/B VGND VGND VPWR VPWR _15362_/X sky130_fd_sc_hd__or4_4
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _25405_/Q VGND VGND VPWR VPWR _12683_/A sky130_fd_sc_hd__inv_2
XFILLER_129_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21846__A2 _13496_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17101_ _17033_/C _17100_/X VGND VGND VPWR VPWR _17105_/B sky130_fd_sc_hd__or2_4
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313_ _25163_/Q _14302_/X _25162_/Q _14307_/X VGND VGND VPWR VPWR _14313_/X sky130_fd_sc_hd__o22a_4
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18081_ _17999_/A _19047_/A VGND VGND VPWR VPWR _18082_/C sky130_fd_sc_hd__or2_4
XANTENNA__18397__A1_N _16223_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15293_ _24991_/Q VGND VGND VPWR VPWR _15309_/A sky130_fd_sc_hd__inv_2
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12905__A _12849_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17032_ _24374_/Q VGND VGND VPWR VPWR _17033_/D sky130_fd_sc_hd__inv_2
X_14244_ _13952_/A _13913_/Y _13893_/B _14244_/D VGND VGND VPWR VPWR _14244_/X sky130_fd_sc_hd__and4_4
XANTENNA__24437__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14175_ _14169_/Y _14110_/X _14111_/X _14174_/X VGND VGND VPWR VPWR _14176_/A sky130_fd_sc_hd__o22a_4
XANTENNA__19672__B1 _19547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13126_ _13126_/A _13126_/B VGND VGND VPWR VPWR _13127_/B sky130_fd_sc_hd__or2_4
XFILLER_125_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18983_ _18982_/Y _18978_/X _18940_/X _18978_/X VGND VGND VPWR VPWR _23886_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24090__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13057_ _13057_/A _13067_/B VGND VGND VPWR VPWR _13064_/B sky130_fd_sc_hd__or2_4
X_17934_ _17930_/A _23884_/Q VGND VGND VPWR VPWR _17934_/X sky130_fd_sc_hd__or2_4
XFILLER_87_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12008_ _11994_/B VGND VGND VPWR VPWR _12008_/Y sky130_fd_sc_hd__inv_2
X_17865_ _17865_/A VGND VGND VPWR VPWR _17865_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21782__A1 _21816_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19604_ _23670_/Q VGND VGND VPWR VPWR _19604_/Y sky130_fd_sc_hd__inv_2
X_16816_ _16807_/A VGND VGND VPWR VPWR _16816_/X sky130_fd_sc_hd__buf_2
X_17796_ _17742_/A _17795_/Y VGND VGND VPWR VPWR _17796_/X sky130_fd_sc_hd__or2_4
XFILLER_94_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25296__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19535_ _13595_/A _14192_/A VGND VGND VPWR VPWR _19535_/X sky130_fd_sc_hd__or2_4
X_13959_ _13958_/X VGND VGND VPWR VPWR _13959_/Y sky130_fd_sc_hd__inv_2
X_16747_ _24455_/Q VGND VGND VPWR VPWR _16747_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21534__A1 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25225__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21534__B2 _21533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18039__A _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16678_ _24483_/Q VGND VGND VPWR VPWR _16678_/Y sky130_fd_sc_hd__inv_2
X_19466_ _19466_/A VGND VGND VPWR VPWR _22339_/B sky130_fd_sc_hd__inv_2
XFILLER_61_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22784__A _22913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18417_ _24643_/Q _18416_/A _16246_/Y _18416_/Y VGND VGND VPWR VPWR _18417_/X sky130_fd_sc_hd__o22a_4
X_15629_ _15629_/A VGND VGND VPWR VPWR _15629_/Y sky130_fd_sc_hd__inv_2
X_19397_ _19396_/Y _19392_/X _19307_/X _19384_/A VGND VGND VPWR VPWR _19397_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16782__A _16781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18348_ _24188_/Q VGND VGND VPWR VPWR _18348_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11786__B1 _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18279_ _24205_/Q VGND VGND VPWR VPWR _18280_/A sky130_fd_sc_hd__inv_2
XANTENNA__12312__A2_N _24807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20310_ _20310_/A VGND VGND VPWR VPWR _20310_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24860__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14724__B1 _21643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21290_ _21302_/A _21289_/X _21290_/C VGND VGND VPWR VPWR _21290_/X sky130_fd_sc_hd__and3_4
XANTENNA__24178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20241_ _20240_/Y _20238_/X _15766_/X _20238_/X VGND VGND VPWR VPWR _23441_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22262__A2 _22224_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18502__A _24172_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16477__B1 _16300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20172_ _23467_/Q VGND VGND VPWR VPWR _20172_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24980_ _24980_/CLK _24980_/D HRESETn VGND VGND VPWR VPWR _24980_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_130_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16229__B1 _16228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23931_ _25205_/CLK _23931_/D HRESETn VGND VGND VPWR VPWR _20537_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15861__A _21026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21582__B _21582_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23862_ _25488_/CLK _23862_/D VGND VGND VPWR VPWR _23862_/Q sky130_fd_sc_hd__dfxtp_4
X_22813_ _24519_/Q _22523_/X _22524_/X _22812_/X VGND VGND VPWR VPWR _22814_/C sky130_fd_sc_hd__a211o_4
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23793_ _24396_/CLK _23793_/D VGND VGND VPWR VPWR _23793_/Q sky130_fd_sc_hd__dfxtp_4
X_25532_ _24691_/CLK _11765_/X HRESETn VGND VGND VPWR VPWR _11763_/A sky130_fd_sc_hd__dfrtp_4
X_22744_ _21064_/A _22741_/X _22705_/A _22743_/X VGND VGND VPWR VPWR _22744_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_53_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_142_0_HCLK clkbuf_7_71_0_HCLK/X VGND VGND VPWR VPWR _23635_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_41_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25463_ _24373_/CLK _25463_/D HRESETn VGND VGND VPWR VPWR _25463_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_94_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22675_ _22674_/X VGND VGND VPWR VPWR _22675_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24948__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24414_ _24413_/CLK _16833_/X HRESETn VGND VGND VPWR VPWR _16832_/A sky130_fd_sc_hd__dfrtp_4
X_21626_ _21596_/A _21626_/B VGND VGND VPWR VPWR _21628_/B sky130_fd_sc_hd__or2_4
XFILLER_90_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21828__A2 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25394_ _25397_/CLK _25394_/D HRESETn VGND VGND VPWR VPWR _12595_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14924__B _14917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21103__A _21103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24345_ _24345_/CLK _24345_/D HRESETn VGND VGND VPWR VPWR _22815_/A sky130_fd_sc_hd__dfrtp_4
X_21557_ _16263_/Y _16449_/A _15115_/A _16723_/A VGND VGND VPWR VPWR _21558_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_14_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20508_ _20506_/X _20507_/X _20602_/A VGND VGND VPWR VPWR _20508_/X sky130_fd_sc_hd__o21a_4
X_12290_ _12290_/A _12290_/B VGND VGND VPWR VPWR _12290_/X sky130_fd_sc_hd__or2_4
X_24276_ _24275_/CLK _24276_/D HRESETn VGND VGND VPWR VPWR _23314_/A sky130_fd_sc_hd__dfrtp_4
X_21488_ _21648_/A _19631_/Y VGND VGND VPWR VPWR _21489_/C sky130_fd_sc_hd__or2_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24530__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23227_ _15567_/Y _22872_/B VGND VGND VPWR VPWR _23227_/X sky130_fd_sc_hd__and2_4
X_20439_ _23922_/Q VGND VGND VPWR VPWR _20439_/X sky130_fd_sc_hd__buf_2
XANTENNA__23312__A1_N _22534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19654__B1 _19553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16468__B1 _16380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12741__A2 _12394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21461__B1 _17722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23158_ _23156_/X _23158_/B _23117_/C VGND VGND VPWR VPWR _23158_/X sky130_fd_sc_hd__or3_4
XFILLER_84_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22109_ _21560_/X _22107_/X _21566_/X _22108_/X VGND VGND VPWR VPWR _22109_/X sky130_fd_sc_hd__o22a_4
X_15980_ _12210_/Y _15978_/X _15620_/X _15978_/X VGND VGND VPWR VPWR _15980_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23202__A1 _24529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12460__A _12235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23089_ _12772_/Y _22707_/X _22272_/X _12539_/Y _22844_/X VGND VGND VPWR VPWR _23089_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14931_ _15179_/A _14930_/A _15180_/A _14930_/Y VGND VGND VPWR VPWR _14939_/B sky130_fd_sc_hd__o22a_4
XFILLER_102_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14862_ _14828_/X _14861_/X _15470_/A _14831_/A VGND VGND VPWR VPWR _14862_/Y sky130_fd_sc_hd__a22oi_4
X_17650_ _17567_/D _17626_/B _17601_/X _17648_/B VGND VGND VPWR VPWR _17651_/A sky130_fd_sc_hd__a211o_4
XANTENNA__19243__A _19242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13813_ _13813_/A _13813_/B VGND VGND VPWR VPWR _15851_/B sky130_fd_sc_hd__or2_4
X_16601_ _16583_/A VGND VGND VPWR VPWR _16601_/X sky130_fd_sc_hd__buf_2
X_17581_ _17569_/X _17611_/B VGND VGND VPWR VPWR _17581_/X sky130_fd_sc_hd__or2_4
X_14793_ _14792_/X VGND VGND VPWR VPWR _14793_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22713__B1 _11802_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16532_ _16530_/Y _16524_/X _16355_/X _16531_/X VGND VGND VPWR VPWR _16532_/X sky130_fd_sc_hd__a2bb2o_4
X_19320_ _18066_/B VGND VGND VPWR VPWR _19320_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11804__A _11803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13744_ _13744_/A _13744_/B _16173_/B _13588_/X VGND VGND VPWR VPWR _14705_/A sky130_fd_sc_hd__or4_4
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16463_ _24564_/Q VGND VGND VPWR VPWR _16463_/Y sky130_fd_sc_hd__inv_2
X_19251_ _23793_/Q VGND VGND VPWR VPWR _19251_/Y sky130_fd_sc_hd__inv_2
X_13675_ _13536_/Y _23343_/B _25285_/Q VGND VGND VPWR VPWR _13675_/X sky130_fd_sc_hd__a21o_4
XANTENNA__15746__A2 _15742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15414_ _15388_/C _15421_/A VGND VGND VPWR VPWR _15423_/A sky130_fd_sc_hd__or2_4
X_18202_ _18202_/A _18198_/X _18201_/X VGND VGND VPWR VPWR _18210_/B sky130_fd_sc_hd__or3_4
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24689__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12626_ _12512_/Y _12626_/B VGND VGND VPWR VPWR _12626_/X sky130_fd_sc_hd__or2_4
X_19182_ _19180_/Y _19176_/X _19136_/X _19181_/X VGND VGND VPWR VPWR _23818_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16394_ _16389_/A VGND VGND VPWR VPWR _16394_/X sky130_fd_sc_hd__buf_2
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18133_ _18133_/A _18133_/B VGND VGND VPWR VPWR _18134_/C sky130_fd_sc_hd__or2_4
XANTENNA__24618__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15345_ _24986_/Q _15345_/B VGND VGND VPWR VPWR _15345_/X sky130_fd_sc_hd__or2_4
XFILLER_40_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12557_ _12557_/A _12557_/B _12557_/C _12557_/D VGND VGND VPWR VPWR _12558_/D sky130_fd_sc_hd__or4_4
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18064_ _18133_/A _23745_/Q VGND VGND VPWR VPWR _18064_/X sky130_fd_sc_hd__or2_4
X_15276_ _15276_/A VGND VGND VPWR VPWR _24999_/D sky130_fd_sc_hd__inv_2
XFILLER_8_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21948__A _21681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12488_ _12269_/Y _12491_/B VGND VGND VPWR VPWR _12492_/B sky130_fd_sc_hd__or2_4
X_17015_ _16059_/Y _16960_/A _16069_/Y _17039_/A VGND VGND VPWR VPWR _17016_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24271__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14227_ _14226_/Y _14224_/X _13837_/X _14224_/X VGND VGND VPWR VPWR _14227_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24200__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14158_ _14144_/X _14157_/Y _14100_/A _14144_/X VGND VGND VPWR VPWR _25203_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13109_ _12993_/A _13107_/X VGND VGND VPWR VPWR _13110_/B sky130_fd_sc_hd__or2_4
X_14089_ _14081_/A VGND VGND VPWR VPWR _14089_/X sky130_fd_sc_hd__buf_2
X_18966_ _18965_/Y _18960_/X _17443_/X _18946_/Y VGND VGND VPWR VPWR _23893_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25477__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17917_ _17911_/Y _13541_/X _17914_/Y _17911_/A _17916_/X VGND VGND VPWR VPWR _24240_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_26_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18897_ _18897_/A VGND VGND VPWR VPWR _22363_/B sky130_fd_sc_hd__inv_2
XFILLER_78_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25406__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17848_ _17750_/D _17848_/B VGND VGND VPWR VPWR _17848_/X sky130_fd_sc_hd__or2_4
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20299__A _20298_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17779_ _17738_/X _17779_/B _17779_/C VGND VGND VPWR VPWR _24274_/D sky130_fd_sc_hd__and3_4
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22704__B1 _21103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18992__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11714__A _24061_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19518_ _23699_/Q VGND VGND VPWR VPWR _22227_/B sky130_fd_sc_hd__inv_2
XFILLER_35_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20790_ _20790_/A VGND VGND VPWR VPWR _20790_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19449_ _17989_/B VGND VGND VPWR VPWR _19449_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_215_0_HCLK clkbuf_8_215_0_HCLK/A VGND VGND VPWR VPWR _24995_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__17401__A _17401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22460_ _20713_/A _21587_/X _15616_/Y _22442_/X VGND VGND VPWR VPWR _22460_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24359__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21411_ _23100_/A VGND VGND VPWR VPWR _22287_/A sky130_fd_sc_hd__buf_2
X_22391_ _22384_/Y _22389_/X _22390_/X _24220_/Q _18235_/A VGND VGND VPWR VPWR _22391_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16017__A _24726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22961__B _22942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16698__B1 _16600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24130_ _24555_/CLK _18762_/X HRESETn VGND VGND VPWR VPWR _24130_/Q sky130_fd_sc_hd__dfrtp_4
X_21342_ _21341_/X VGND VGND VPWR VPWR _21343_/D sky130_fd_sc_hd__inv_2
XFILLER_120_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18857__A1_N _16503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24061_ _23370_/CLK _24061_/D HRESETn VGND VGND VPWR VPWR _24061_/Q sky130_fd_sc_hd__dfrtp_4
X_21273_ _21273_/A VGND VGND VPWR VPWR _21273_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23012_ _12886_/A _21872_/X _16943_/Y _22821_/X VGND VGND VPWR VPWR _23012_/X sky130_fd_sc_hd__o22a_4
X_20224_ _20211_/Y VGND VGND VPWR VPWR _20224_/X sky130_fd_sc_hd__buf_2
XFILLER_103_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20797__A2 _20676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20155_ _22075_/B _20149_/X _20085_/X _20154_/X VGND VGND VPWR VPWR _23474_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14910__D _14909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23994__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23923__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20086_ _20095_/A VGND VGND VPWR VPWR _20086_/X sky130_fd_sc_hd__buf_2
X_24963_ _24977_/CLK _15425_/Y HRESETn VGND VGND VPWR VPWR _24963_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25147__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12430__D _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19063__A _19062_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23914_ _23434_/CLK _23914_/D VGND VGND VPWR VPWR _18906_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24894_ _24909_/CLK _15603_/X HRESETn VGND VGND VPWR VPWR _24894_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23845_ _23847_/CLK _19103_/X VGND VGND VPWR VPWR _23845_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20002__A _20014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12239__B2 _24749_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_25_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_11790_ _25524_/Q VGND VGND VPWR VPWR _11790_/Y sky130_fd_sc_hd__inv_2
X_23776_ _23618_/CLK _19300_/X VGND VGND VPWR VPWR _19299_/A sky130_fd_sc_hd__dfxtp_4
X_20988_ scl_oen_o_S5 _20988_/B VGND VGND VPWR VPWR _20988_/X sky130_fd_sc_hd__and2_4
XFILLER_53_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25515_ _25514_/CLK _11830_/X HRESETn VGND VGND VPWR VPWR _11828_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_13_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23313__A _23281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22727_ _11664_/Y _22727_/B VGND VGND VPWR VPWR _22727_/X sky130_fd_sc_hd__and2_4
XANTENNA__24782__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13460_ _13428_/A _13458_/X _13459_/X VGND VGND VPWR VPWR _13460_/X sky130_fd_sc_hd__and3_4
X_25446_ _25449_/CLK _12413_/Y HRESETn VGND VGND VPWR VPWR _12191_/A sky130_fd_sc_hd__dfrtp_4
X_22658_ _22658_/A _22658_/B _22649_/X _22658_/D VGND VGND VPWR VPWR _22658_/X sky130_fd_sc_hd__or4_4
X_12411_ _12290_/B _12391_/B _12290_/A VGND VGND VPWR VPWR _12411_/X sky130_fd_sc_hd__o21a_4
XFILLER_51_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24711__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21609_ _21609_/A _21607_/X _21608_/X VGND VGND VPWR VPWR _21609_/X sky130_fd_sc_hd__and3_4
X_13391_ _13455_/A _19719_/A VGND VGND VPWR VPWR _13393_/B sky130_fd_sc_hd__or2_4
X_25377_ _25368_/CLK _12900_/Y HRESETn VGND VGND VPWR VPWR _25377_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12455__A _12249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22589_ _22549_/A _22589_/B VGND VGND VPWR VPWR _22589_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24029__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15130_ _24977_/Q VGND VGND VPWR VPWR _15130_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16689__B1 _15747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12342_ _13102_/A VGND VGND VPWR VPWR _12995_/A sky130_fd_sc_hd__inv_2
XFILLER_51_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21682__B1 _21493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24328_ _24330_/CLK _24328_/D HRESETn VGND VGND VPWR VPWR _17242_/A sky130_fd_sc_hd__dfrtp_4
X_15061_ _14885_/Y _14942_/Y _15249_/A _15061_/D VGND VGND VPWR VPWR _15064_/C sky130_fd_sc_hd__or4_4
XANTENNA__15766__A _15766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12273_ _12273_/A _12273_/B VGND VGND VPWR VPWR _12390_/B sky130_fd_sc_hd__or2_4
X_24259_ _24682_/CLK _24259_/D HRESETn VGND VGND VPWR VPWR _24259_/Q sky130_fd_sc_hd__dfrtp_4
X_14012_ _14012_/A _14007_/X _14012_/C _14040_/C VGND VGND VPWR VPWR _14012_/X sky130_fd_sc_hd__or4_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12902__B _12799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18820_ _18742_/A _18820_/B _18819_/Y VGND VGND VPWR VPWR _18820_/X sky130_fd_sc_hd__and3_4
XANTENNA__17981__A _18087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12190__A _22550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18751_ _18656_/Y _18745_/X _18733_/X _18747_/Y VGND VGND VPWR VPWR _18752_/A sky130_fd_sc_hd__a211o_4
XANTENNA__12478__A1 _12282_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15963_ _12200_/Y _15960_/X _15962_/X _15960_/X VGND VGND VPWR VPWR _15963_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_107_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_215_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16597__A _16597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17702_ _17702_/A VGND VGND VPWR VPWR _17735_/B sky130_fd_sc_hd__inv_2
X_14914_ _25013_/Q _14913_/A _15219_/A _14913_/Y VGND VGND VPWR VPWR _14924_/A sky130_fd_sc_hd__o22a_4
XFILLER_64_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15894_ _15894_/A VGND VGND VPWR VPWR _15894_/X sky130_fd_sc_hd__buf_2
X_18682_ _18682_/A _18682_/B _18639_/Y VGND VGND VPWR VPWR _18683_/D sky130_fd_sc_hd__or3_4
XFILLER_110_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22111__B _22111_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17633_ _17633_/A VGND VGND VPWR VPWR _17633_/Y sky130_fd_sc_hd__inv_2
X_14845_ _14831_/A VGND VGND VPWR VPWR _14845_/X sky130_fd_sc_hd__buf_2
XFILLER_63_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14776_ _25045_/Q _14776_/B VGND VGND VPWR VPWR _14783_/A sky130_fd_sc_hd__and2_4
X_17564_ _24294_/Q VGND VGND VPWR VPWR _17564_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11988_ _11654_/B _11977_/X _11987_/Y VGND VGND VPWR VPWR _11988_/X sky130_fd_sc_hd__o21a_4
X_19303_ _19301_/Y _19302_/X _19212_/X _19302_/X VGND VGND VPWR VPWR _19303_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22162__B2 _14220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13727_ _11669_/Y _13683_/B VGND VGND VPWR VPWR _13727_/Y sky130_fd_sc_hd__nand2_4
X_16515_ _24543_/Q VGND VGND VPWR VPWR _16515_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17495_ _25513_/Q _17494_/Y _11756_/Y _17605_/A VGND VGND VPWR VPWR _17495_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19234_ _13372_/B VGND VGND VPWR VPWR _19234_/Y sky130_fd_sc_hd__inv_2
X_13658_ _13658_/A _13658_/B VGND VGND VPWR VPWR _13659_/B sky130_fd_sc_hd__or2_4
X_16446_ _16445_/Y _16375_/A _16366_/X _16375_/A VGND VGND VPWR VPWR _24567_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24452__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12609_ _12609_/A _12679_/A _12576_/Y _12567_/Y VGND VGND VPWR VPWR _12609_/X sky130_fd_sc_hd__or4_4
XFILLER_73_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16377_ _16368_/Y _16375_/X _16376_/X _16375_/X VGND VGND VPWR VPWR _24598_/D sky130_fd_sc_hd__a2bb2o_4
X_19165_ _19164_/Y _19160_/X _19117_/X _19160_/X VGND VGND VPWR VPWR _23824_/D sky130_fd_sc_hd__a2bb2o_4
X_13589_ _13588_/X VGND VGND VPWR VPWR _14555_/B sky130_fd_sc_hd__inv_2
Xclkbuf_8_45_0_HCLK clkbuf_8_45_0_HCLK/A VGND VGND VPWR VPWR _23689_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15328_ _15310_/B _15308_/X VGND VGND VPWR VPWR _15329_/A sky130_fd_sc_hd__or2_4
X_18116_ _17999_/A _19049_/A VGND VGND VPWR VPWR _18117_/C sky130_fd_sc_hd__or2_4
XFILLER_8_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19096_ _21753_/B _19091_/X _16881_/X _19091_/X VGND VGND VPWR VPWR _23848_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15259_ _15251_/B _15250_/X VGND VGND VPWR VPWR _15262_/B sky130_fd_sc_hd__or2_4
X_18047_ _18005_/A _18045_/X _18047_/C VGND VGND VPWR VPWR _18048_/C sky130_fd_sc_hd__and3_4
XFILLER_67_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24945__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13196__A _13195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21976__B2 _20331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11709__A _11707_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18841__A1 _24564_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19998_ _19997_/Y _19991_/X _19885_/X _19991_/A VGND VGND VPWR VPWR _23533_/D sky130_fd_sc_hd__a2bb2o_4
X_18949_ _13222_/B VGND VGND VPWR VPWR _18949_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25240__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21960_ _21957_/X _21958_/X _21959_/X VGND VGND VPWR VPWR _21960_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_132_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16300__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20911_ _24050_/Q _24049_/Q _20889_/B _20900_/B VGND VGND VPWR VPWR _20911_/X sky130_fd_sc_hd__or4_4
X_21891_ _21886_/A _18909_/Y VGND VGND VPWR VPWR _21891_/X sky130_fd_sc_hd__or2_4
XFILLER_55_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18609__A2_N _18608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23630_ _23388_/CLK _23630_/D VGND VGND VPWR VPWR _23630_/Q sky130_fd_sc_hd__dfxtp_4
X_20842_ _13658_/A _13658_/B _20852_/B VGND VGND VPWR VPWR _20842_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_81_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23561_ _25264_/CLK _19919_/X VGND VGND VPWR VPWR _19918_/A sky130_fd_sc_hd__dfxtp_4
X_20773_ _20771_/Y _20767_/X _20772_/X VGND VGND VPWR VPWR _20773_/X sky130_fd_sc_hd__o21a_4
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25300_ _25301_/CLK _25300_/D HRESETn VGND VGND VPWR VPWR _25300_/Q sky130_fd_sc_hd__dfrtp_4
X_22512_ _16697_/Y _21428_/X VGND VGND VPWR VPWR _22512_/X sky130_fd_sc_hd__and2_4
XFILLER_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23492_ _23434_/CLK _20107_/X VGND VGND VPWR VPWR _20103_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22972__A _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24193__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25231_ _24151_/CLK _25231_/D HRESETn VGND VGND VPWR VPWR _21142_/A sky130_fd_sc_hd__dfrtp_4
X_22443_ _15008_/Y _21067_/X _16728_/A _14916_/Y _22442_/X VGND VGND VPWR VPWR _22443_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__15591__B1 _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19857__B1 _19790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24122__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21588__A _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25162_ _25305_/CLK _25162_/D HRESETn VGND VGND VPWR VPWR _25162_/Q sky130_fd_sc_hd__dfrtp_4
X_22374_ _22050_/X _20146_/Y VGND VGND VPWR VPWR _22374_/X sky130_fd_sc_hd__or2_4
X_24113_ _24120_/CLK _24113_/D HRESETn VGND VGND VPWR VPWR _18679_/A sky130_fd_sc_hd__dfrtp_4
X_21325_ _21325_/A VGND VGND VPWR VPWR _22798_/A sky130_fd_sc_hd__buf_2
XANTENNA__14490__A _25102_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25093_ _25093_/CLK _14525_/X HRESETn VGND VGND VPWR VPWR _21841_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25399__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24044_ _24496_/CLK _24044_/D HRESETn VGND VGND VPWR VPWR _24044_/Q sky130_fd_sc_hd__dfrtp_4
X_21256_ _21253_/A _21256_/B VGND VGND VPWR VPWR _21257_/C sky130_fd_sc_hd__or2_4
XFILLER_89_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25328__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20207_ _23453_/Q VGND VGND VPWR VPWR _21231_/B sky130_fd_sc_hd__inv_2
XFILLER_81_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21187_ _21183_/X _21186_/X _17720_/X VGND VGND VPWR VPWR _21196_/B sky130_fd_sc_hd__o21a_4
XFILLER_132_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16843__B1 _16521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20138_ _21772_/B _20133_/X _20092_/X _20133_/X VGND VGND VPWR VPWR _23480_/D sky130_fd_sc_hd__a2bb2o_4
X_12960_ _12833_/Y _12960_/B VGND VGND VPWR VPWR _12964_/B sky130_fd_sc_hd__or2_4
X_20069_ _20064_/X _18326_/X _11842_/A _13273_/B _20066_/X VGND VGND VPWR VPWR _23506_/D
+ sky130_fd_sc_hd__a32o_4
X_24946_ _24950_/CLK _15460_/X HRESETn VGND VGND VPWR VPWR _13927_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_38_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11911_ _11910_/X VGND VGND VPWR VPWR _11916_/B sky130_fd_sc_hd__inv_2
XFILLER_46_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18060__A2 _18040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12891_ _12749_/Y _12889_/A VGND VGND VPWR VPWR _12891_/X sky130_fd_sc_hd__or2_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24877_ _24909_/CLK _24877_/D HRESETn VGND VGND VPWR VPWR _24877_/Q sky130_fd_sc_hd__dfrtp_4
X_14630_ _14614_/X _14630_/B VGND VGND VPWR VPWR _14630_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24963__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11842_ _11842_/A VGND VGND VPWR VPWR _11842_/X sky130_fd_sc_hd__buf_2
XFILLER_79_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19521__A _19528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23828_ _23828_/CLK _23828_/D VGND VGND VPWR VPWR _23828_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24064__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14561_ _14561_/A _14560_/X VGND VGND VPWR VPWR _14561_/X sky130_fd_sc_hd__or2_4
XFILLER_14_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11773_ _25529_/Q VGND VGND VPWR VPWR _11773_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20155__B1 _20085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23759_ _23722_/CLK _23759_/D VGND VGND VPWR VPWR _18150_/B sky130_fd_sc_hd__dfxtp_4
X_13512_ _13497_/Y VGND VGND VPWR VPWR _13512_/X sky130_fd_sc_hd__buf_2
X_16300_ HWDATA[25] VGND VGND VPWR VPWR _16300_/X sky130_fd_sc_hd__buf_2
X_17280_ _17261_/B _17269_/C _17279_/X _17276_/B VGND VGND VPWR VPWR _17280_/X sky130_fd_sc_hd__a211o_4
XFILLER_92_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14492_ _25101_/Q VGND VGND VPWR VPWR _14492_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16231_ _11803_/X VGND VGND VPWR VPWR _16231_/X sky130_fd_sc_hd__buf_2
XFILLER_110_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13443_ _13379_/A _23901_/Q VGND VGND VPWR VPWR _13443_/X sky130_fd_sc_hd__or2_4
X_25429_ _25449_/CLK _25429_/D HRESETn VGND VGND VPWR VPWR _25429_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15582__B1 _11771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19848__B1 _19777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17976__A _17990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16880__A _16880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_4_0_HCLK clkbuf_8_5_0_HCLK/A VGND VGND VPWR VPWR _23847_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16162_ _16161_/Y _16157_/X _15986_/X _16157_/X VGND VGND VPWR VPWR _24670_/D sky130_fd_sc_hd__a2bb2o_4
X_13374_ _13301_/X _13372_/X _13374_/C VGND VGND VPWR VPWR _13374_/X sky130_fd_sc_hd__and3_4
XFILLER_16_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15113_ _15111_/A _24576_/Q _15299_/A _15112_/Y VGND VGND VPWR VPWR _15113_/X sky130_fd_sc_hd__o22a_4
X_12325_ _25329_/Q _24814_/Q _13096_/A _12324_/Y VGND VGND VPWR VPWR _12325_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16093_ _16087_/A VGND VGND VPWR VPWR _16094_/A sky130_fd_sc_hd__buf_2
XFILLER_126_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15044_ _14949_/Y VGND VGND VPWR VPWR _15210_/B sky130_fd_sc_hd__buf_2
X_19921_ _19920_/Y _19916_/X _19790_/X _19916_/X VGND VGND VPWR VPWR _19921_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12256_ _12278_/C _24739_/Q _25448_/Q _12255_/Y VGND VGND VPWR VPWR _12262_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12699__A1 _12565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25069__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19852_ _19859_/A VGND VGND VPWR VPWR _19852_/X sky130_fd_sc_hd__buf_2
X_12187_ _12187_/A VGND VGND VPWR VPWR _12188_/A sky130_fd_sc_hd__inv_2
X_18803_ _18782_/X _18803_/B VGND VGND VPWR VPWR _18803_/X sky130_fd_sc_hd__or2_4
X_19783_ _16872_/A VGND VGND VPWR VPWR _19783_/X sky130_fd_sc_hd__buf_2
XFILLER_122_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16995_ _24704_/Q _16993_/Y _24708_/Q _17130_/A VGND VGND VPWR VPWR _16998_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18734_ _18675_/X _18728_/B _18733_/X _18729_/Y VGND VGND VPWR VPWR _18734_/X sky130_fd_sc_hd__a211o_4
XFILLER_95_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15946_ _12194_/Y _15939_/X _15944_/X _15945_/X VGND VGND VPWR VPWR _15946_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18665_ _16608_/Y _18601_/A _16616_/Y _18681_/A VGND VGND VPWR VPWR _18665_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15877_ _15850_/X _15857_/X _15729_/X _24795_/Q _15864_/X VGND VGND VPWR VPWR _24795_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17616_ _17616_/A _17616_/B VGND VGND VPWR VPWR _17617_/C sky130_fd_sc_hd__nand2_4
X_14828_ _14810_/A VGND VGND VPWR VPWR _14828_/X sky130_fd_sc_hd__buf_2
X_18596_ _18595_/X VGND VGND VPWR VPWR _18596_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16584__A1_N _16581_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24633__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17547_ _11745_/Y _24308_/Q _11745_/Y _24308_/Q VGND VGND VPWR VPWR _17550_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14759_ _21608_/A _14746_/B _14752_/X VGND VGND VPWR VPWR _14759_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_32_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17478_ _17477_/Y VGND VGND VPWR VPWR _17478_/X sky130_fd_sc_hd__buf_2
XANTENNA__22792__A _22792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19217_ _19216_/Y _19211_/X _19149_/X _19197_/X VGND VGND VPWR VPWR _19217_/X sky130_fd_sc_hd__a2bb2o_4
X_16429_ _16433_/A VGND VGND VPWR VPWR _16429_/X sky130_fd_sc_hd__buf_2
XANTENNA__15573__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19839__B1 _19797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16790__A _24434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21646__B1 _13784_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19148_ _23829_/Q VGND VGND VPWR VPWR _19148_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18511__B1 _18487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19079_ _13401_/B VGND VGND VPWR VPWR _19079_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25492__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21110_ _21030_/X _21109_/X _13141_/Y _15665_/A VGND VGND VPWR VPWR _21110_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22090_ _22923_/A VGND VGND VPWR VPWR _22090_/X sky130_fd_sc_hd__buf_2
XFILLER_133_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25421__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21041_ _24842_/Q _21021_/X _21024_/X _21040_/X VGND VGND VPWR VPWR _21042_/C sky130_fd_sc_hd__a211o_4
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18510__A _18460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12236__A1_N _12235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24800_ _24800_/CLK _15871_/X HRESETn VGND VGND VPWR VPWR _23213_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_68_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22992_ _22992_/A _22796_/B VGND VGND VPWR VPWR _22995_/B sky130_fd_sc_hd__or2_4
X_24731_ _24355_/CLK _16006_/X HRESETn VGND VGND VPWR VPWR _24731_/Q sky130_fd_sc_hd__dfrtp_4
X_21943_ _21454_/A _21941_/X _21942_/X VGND VGND VPWR VPWR _21943_/X sky130_fd_sc_hd__and3_4
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22982__A1_N _17252_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_7_0_HCLK_A clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24662_ _24162_/CLK _24662_/D HRESETn VGND VGND VPWR VPWR _23232_/A sky130_fd_sc_hd__dfrtp_4
X_21874_ _25424_/Q _23271_/A _21873_/X _21095_/X VGND VGND VPWR VPWR _21874_/X sky130_fd_sc_hd__a211o_4
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24374__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _23598_/CLK _19772_/X VGND VGND VPWR VPWR _13458_/B sky130_fd_sc_hd__dfxtp_4
X_20825_ _13653_/A _13653_/B _13655_/B VGND VGND VPWR VPWR _20825_/X sky130_fd_sc_hd__o21a_4
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24593_ _24995_/CLK _16390_/X HRESETn VGND VGND VPWR VPWR _24593_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13811__B1 _13810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17002__B1 _16037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24303__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11902__A RsRx_S1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23544_ _23533_/CLK _23544_/D VGND VGND VPWR VPWR _23544_/Q sky130_fd_sc_hd__dfxtp_4
X_20756_ _20743_/X _20755_/Y _15595_/A _20747_/X VGND VGND VPWR VPWR _24014_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15564__B1 _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23475_ _23467_/CLK _23475_/D VGND VGND VPWR VPWR _23475_/Q sky130_fd_sc_hd__dfxtp_4
X_20687_ _13121_/Y _13123_/B _13124_/Y VGND VGND VPWR VPWR _20687_/X sky130_fd_sc_hd__o21a_4
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25214_ _24322_/CLK _25214_/D HRESETn VGND VGND VPWR VPWR _14003_/C sky130_fd_sc_hd__dfrtp_4
X_22426_ _21312_/X VGND VGND VPWR VPWR _22426_/X sky130_fd_sc_hd__buf_2
XFILLER_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15731__A1_N _12586_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25509__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25145_ _25141_/CLK _25145_/D HRESETn VGND VGND VPWR VPWR _25145_/Q sky130_fd_sc_hd__dfrtp_4
X_22357_ _22068_/A _22357_/B VGND VGND VPWR VPWR _22357_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_91_0_HCLK clkbuf_8_91_0_HCLK/A VGND VGND VPWR VPWR _24502_/CLK sky130_fd_sc_hd__clkbuf_1
X_12110_ _12109_/Y _12107_/X _11838_/X _12107_/X VGND VGND VPWR VPWR _12110_/X sky130_fd_sc_hd__a2bb2o_4
X_21308_ _21275_/X _21286_/X _21290_/X _21301_/X _21307_/X VGND VGND VPWR VPWR _21510_/A
+ sky130_fd_sc_hd__o41a_4
X_13090_ _12992_/Y _13086_/X VGND VGND VPWR VPWR _13090_/Y sky130_fd_sc_hd__nand2_4
X_25076_ _25290_/CLK _14600_/X HRESETn VGND VGND VPWR VPWR _25076_/Q sky130_fd_sc_hd__dfrtp_4
X_22288_ _22764_/A VGND VGND VPWR VPWR _22288_/X sky130_fd_sc_hd__buf_2
XFILLER_2_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22305__A1_N _14381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12041_ _12034_/A VGND VGND VPWR VPWR _12041_/X sky130_fd_sc_hd__buf_2
XFILLER_105_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24027_ _24025_/CLK _20810_/X HRESETn VGND VGND VPWR VPWR _13137_/C sky130_fd_sc_hd__dfrtp_4
X_21239_ _14680_/X _18918_/Y VGND VGND VPWR VPWR _21239_/X sky130_fd_sc_hd__or2_4
XANTENNA__19516__A _19528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20612__A1 _15473_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15800_ _12328_/Y _15799_/X _11749_/X _15799_/X VGND VGND VPWR VPWR _15800_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17036__A _17036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13992_ _14001_/A _13989_/X _14040_/C VGND VGND VPWR VPWR _13992_/X sky130_fd_sc_hd__or3_4
X_16780_ _14991_/Y _16778_/X _16528_/X _16778_/X VGND VGND VPWR VPWR _24438_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14379__B _18895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21781__A _21781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12943_ _12774_/Y _12833_/Y _12959_/A _12959_/B VGND VGND VPWR VPWR _12944_/D sky130_fd_sc_hd__or4_4
X_15731_ _12586_/Y _15721_/X _11774_/X _15721_/X VGND VGND VPWR VPWR _15731_/X sky130_fd_sc_hd__a2bb2o_4
X_24929_ _24930_/CLK _24929_/D HRESETn VGND VGND VPWR VPWR _15503_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_19_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18450_ _18450_/A _18450_/B _18444_/X _18449_/X VGND VGND VPWR VPWR _18451_/B sky130_fd_sc_hd__or4_4
XFILLER_94_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12874_ _12882_/A VGND VGND VPWR VPWR _12874_/X sky130_fd_sc_hd__buf_2
X_15662_ _15662_/A _15662_/B _21027_/A _15662_/D VGND VGND VPWR VPWR _15670_/A sky130_fd_sc_hd__or4_4
XFILLER_34_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17401_ _17401_/A VGND VGND VPWR VPWR _17401_/X sky130_fd_sc_hd__buf_2
XANTENNA__20391__A3 _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11825_ HWDATA[9] VGND VGND VPWR VPWR _11825_/X sky130_fd_sc_hd__buf_2
X_14613_ _14613_/A VGND VGND VPWR VPWR _14613_/Y sky130_fd_sc_hd__inv_2
X_15593_ _15588_/A VGND VGND VPWR VPWR _15593_/X sky130_fd_sc_hd__buf_2
X_18381_ _18381_/A VGND VGND VPWR VPWR _18381_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14395__A _15986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22668__A2 _22665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11812__A HWDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24044__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14010_/X VGND VGND VPWR VPWR _14545_/C sky130_fd_sc_hd__inv_2
X_17332_ _17252_/A _17330_/A VGND VGND VPWR VPWR _17333_/C sky130_fd_sc_hd__or2_4
XPHY_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11756_/A VGND VGND VPWR VPWR _11756_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _21027_/B _14475_/B VGND VGND VPWR VPWR _14481_/A sky130_fd_sc_hd__nor2_4
X_17263_ _24359_/Q _17263_/B VGND VGND VPWR VPWR _17263_/X sky130_fd_sc_hd__or2_4
XFILLER_109_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _11685_/A _24221_/Q _11685_/Y _11686_/Y VGND VGND VPWR VPWR _11688_/D sky130_fd_sc_hd__o22a_4
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19002_ _23880_/Q VGND VGND VPWR VPWR _19002_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13426_ _13426_/A _13426_/B VGND VGND VPWR VPWR _13426_/X sky130_fd_sc_hd__or2_4
X_16214_ _24654_/Q VGND VGND VPWR VPWR _16214_/Y sky130_fd_sc_hd__inv_2
X_17194_ _23246_/A VGND VGND VPWR VPWR _17194_/Y sky130_fd_sc_hd__inv_2
X_16145_ _16142_/Y _16138_/X _16143_/X _16144_/X VGND VGND VPWR VPWR _16145_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21021__A _22523_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13357_ _13421_/A _13355_/X _13357_/C VGND VGND VPWR VPWR _13357_/X sky130_fd_sc_hd__and3_4
XANTENNA__13739__A _21643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12308_ _12308_/A VGND VGND VPWR VPWR _12308_/Y sky130_fd_sc_hd__inv_2
X_16076_ _16075_/Y _15996_/X _15480_/X _15996_/X VGND VGND VPWR VPWR _16076_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_119_0_HCLK clkbuf_7_59_0_HCLK/X VGND VGND VPWR VPWR _24557_/CLK sky130_fd_sc_hd__clkbuf_1
X_13288_ _13392_/A _13288_/B VGND VGND VPWR VPWR _13288_/X sky130_fd_sc_hd__or2_4
XFILLER_29_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15027_ _15027_/A VGND VGND VPWR VPWR _15027_/Y sky130_fd_sc_hd__inv_2
X_19904_ _23566_/Q VGND VGND VPWR VPWR _19904_/Y sky130_fd_sc_hd__inv_2
X_12239_ _12238_/X _24749_/Q _12238_/A _24749_/Q VGND VGND VPWR VPWR _12239_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19835_ _19835_/A VGND VGND VPWR VPWR _19835_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24885__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19766_ _19751_/Y VGND VGND VPWR VPWR _19766_/X sky130_fd_sc_hd__buf_2
X_16978_ _24367_/Q VGND VGND VPWR VPWR _17038_/C sky130_fd_sc_hd__inv_2
XFILLER_7_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20785__A1_N _20770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18717_ _18772_/A _18695_/X VGND VGND VPWR VPWR _18717_/X sky130_fd_sc_hd__or2_4
XFILLER_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24814__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15929_ _15669_/X _15795_/A _15927_/X _24767_/Q _15928_/X VGND VGND VPWR VPWR _15929_/X
+ sky130_fd_sc_hd__a32o_4
X_19697_ _19697_/A VGND VGND VPWR VPWR _19697_/X sky130_fd_sc_hd__buf_2
XANTENNA__16785__A _16785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18648_ _16565_/Y _18647_/X _16565_/Y _24136_/Q VGND VGND VPWR VPWR _18652_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23305__B1 _24873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20382__A3 _13835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20119__B1 _20096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18579_ _18575_/B _18577_/Y _18582_/C VGND VGND VPWR VPWR _24151_/D sky130_fd_sc_hd__and3_4
XFILLER_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20610_ _17403_/A VGND VGND VPWR VPWR _20611_/C sky130_fd_sc_hd__buf_2
X_21590_ _13653_/A _21588_/X _23999_/Q _21589_/X VGND VGND VPWR VPWR _21590_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17535__B2 _17630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20541_ _20541_/A VGND VGND VPWR VPWR _23932_/D sky130_fd_sc_hd__inv_2
XFILLER_123_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20754__B _20745_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23260_ _22819_/X _23251_/Y _23255_/Y _23259_/X VGND VGND VPWR VPWR _23268_/C sky130_fd_sc_hd__a211o_4
X_20472_ _14205_/A _14207_/A VGND VGND VPWR VPWR _20472_/X sky130_fd_sc_hd__or2_4
XANTENNA__23084__A2 _22833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14752__B _14744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22211_ _14712_/A _22207_/X _22210_/X VGND VGND VPWR VPWR _22211_/X sky130_fd_sc_hd__or3_4
Xclkbuf_7_15_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__22292__B1 _22132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23191_ _12291_/A _22980_/X _17785_/A _22483_/X VGND VGND VPWR VPWR _23191_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_78_0_HCLK clkbuf_7_79_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_78_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15849__A1 _15669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22142_ _21025_/A _22141_/X _22125_/X _12345_/A _15544_/X VGND VGND VPWR VPWR _22142_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_69_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21866__A _11720_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15864__A _15864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22073_ _21763_/A _22071_/X _22072_/X VGND VGND VPWR VPWR _22073_/X sky130_fd_sc_hd__and3_4
XFILLER_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21024_ _21024_/A VGND VGND VPWR VPWR _21024_/X sky130_fd_sc_hd__buf_2
XFILLER_138_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16274__A1 _15655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22697__A _23085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24555__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22975_ _21025_/A VGND VGND VPWR VPWR _22975_/X sky130_fd_sc_hd__buf_2
XANTENNA__16695__A _16645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19071__A _16781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21926_ _21945_/A _21926_/B VGND VGND VPWR VPWR _21926_/X sky130_fd_sc_hd__or2_4
X_24714_ _24318_/CLK _16048_/X HRESETn VGND VGND VPWR VPWR _24714_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24645_ _24643_/CLK _24645_/D HRESETn VGND VGND VPWR VPWR _22583_/A sky130_fd_sc_hd__dfrtp_4
X_21857_ _24571_/Q _23082_/B VGND VGND VPWR VPWR _21861_/B sky130_fd_sc_hd__or2_4
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21307__C1 _21306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12743__A1_N _12842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _20804_/X VGND VGND VPWR VPWR _20808_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23311__A3 _22127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12590_/A VGND VGND VPWR VPWR _12596_/A sky130_fd_sc_hd__inv_2
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24576_ _24572_/CLK _16430_/X HRESETn VGND VGND VPWR VPWR _24576_/Q sky130_fd_sc_hd__dfrtp_4
X_21788_ _21650_/A _21788_/B VGND VGND VPWR VPWR _21788_/X sky130_fd_sc_hd__or2_4
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23527_ _23550_/CLK _20015_/X VGND VGND VPWR VPWR _20013_/A sky130_fd_sc_hd__dfxtp_4
X_20739_ _20740_/B VGND VGND VPWR VPWR _20739_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15537__B1 HADDR[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ _14254_/Y _14259_/X _13835_/X _14259_/X VGND VGND VPWR VPWR _14260_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22807__C1 _22806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23458_ _23609_/CLK _23458_/D VGND VGND VPWR VPWR _23458_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25343__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13211_ _13379_/A _13211_/B VGND VGND VPWR VPWR _13211_/X sky130_fd_sc_hd__or2_4
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22409_ _21741_/A _22409_/B VGND VGND VPWR VPWR _22409_/Y sky130_fd_sc_hd__nor2_4
X_14191_ _13787_/A _19581_/B _11725_/B _13777_/A VGND VGND VPWR VPWR _14192_/A sky130_fd_sc_hd__or4_4
XANTENNA__12463__A _12430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23389_ _23533_/CLK _23389_/D VGND VGND VPWR VPWR _23389_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13142_ _21007_/A _13140_/X _13141_/Y VGND VGND VPWR VPWR _25321_/D sky130_fd_sc_hd__o21a_4
XFILLER_125_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25128_ _25122_/CLK _25128_/D HRESETn VGND VGND VPWR VPWR _25128_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__15774__A _15845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13073_ _13073_/A VGND VGND VPWR VPWR _13073_/Y sky130_fd_sc_hd__inv_2
X_17950_ _14648_/X _17950_/B _17950_/C VGND VGND VPWR VPWR _17950_/X sky130_fd_sc_hd__and3_4
X_25059_ _25044_/CLK _14672_/X HRESETn VGND VGND VPWR VPWR _25059_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_65_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18150__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12024_ _12019_/A _12019_/B _12021_/Y VGND VGND VPWR VPWR _12024_/X sky130_fd_sc_hd__o21a_4
X_16901_ _17785_/A VGND VGND VPWR VPWR _17786_/A sky130_fd_sc_hd__inv_2
X_17881_ _16920_/Y _17878_/B VGND VGND VPWR VPWR _17882_/C sky130_fd_sc_hd__nand2_4
X_19620_ _19617_/Y _19611_/X _19618_/X _19619_/X VGND VGND VPWR VPWR _19620_/X sky130_fd_sc_hd__a2bb2o_4
X_16832_ _16832_/A VGND VGND VPWR VPWR _16832_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14276__B1 _13810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24296__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19551_ _23687_/Q VGND VGND VPWR VPWR _19551_/Y sky130_fd_sc_hd__inv_2
X_16763_ _24447_/Q VGND VGND VPWR VPWR _16763_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13975_ _13975_/A VGND VGND VPWR VPWR _14006_/A sky130_fd_sc_hd__buf_2
XFILLER_93_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22400__A _22400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18502_ _24172_/Q _18506_/B VGND VGND VPWR VPWR _18504_/B sky130_fd_sc_hd__or2_4
XFILLER_74_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24225__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15714_ HWDATA[30] VGND VGND VPWR VPWR _15714_/X sky130_fd_sc_hd__buf_2
XFILLER_47_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12926_ _12926_/A _12926_/B VGND VGND VPWR VPWR _12928_/B sky130_fd_sc_hd__or2_4
X_19482_ _23711_/Q VGND VGND VPWR VPWR _19482_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23215__B _23214_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16694_ _24476_/Q VGND VGND VPWR VPWR _22560_/A sky130_fd_sc_hd__inv_2
XFILLER_62_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18962__B1 _18961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18433_ _16207_/Y _24168_/Q _16207_/Y _24168_/Q VGND VGND VPWR VPWR _18433_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21016__A _21408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15645_ _15648_/A VGND VGND VPWR VPWR _15646_/A sky130_fd_sc_hd__inv_2
X_12857_ _12864_/A _12840_/Y _12830_/Y _12856_/X VGND VGND VPWR VPWR _12858_/A sky130_fd_sc_hd__or4_4
XFILLER_61_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21849__B1 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11808_ HWDATA[13] VGND VGND VPWR VPWR _11809_/A sky130_fd_sc_hd__buf_2
X_18364_ _18356_/X _18363_/Y _24188_/Q _18355_/Y VGND VGND VPWR VPWR _24188_/D sky130_fd_sc_hd__a2bb2o_4
X_12788_ _24774_/Q VGND VGND VPWR VPWR _12788_/Y sky130_fd_sc_hd__inv_2
X_15576_ _15574_/Y _15575_/X _11764_/X _15575_/X VGND VGND VPWR VPWR _15576_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17220_/Y _17309_/X _17279_/X _17311_/Y VGND VGND VPWR VPWR _17315_/X sky130_fd_sc_hd__a211o_4
X_11739_ _11739_/A _22913_/A VGND VGND VPWR VPWR _11739_/X sky130_fd_sc_hd__and2_4
X_14527_ _14521_/X _14526_/X _25104_/Q _14517_/X VGND VGND VPWR VPWR _25092_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15949__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18295_ _18295_/A VGND VGND VPWR VPWR _18295_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17246_ _17196_/Y _17246_/B _17246_/C _17245_/X VGND VGND VPWR VPWR _17247_/D sky130_fd_sc_hd__or4_4
X_14458_ _14458_/A VGND VGND VPWR VPWR _14458_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25084__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13409_ _13345_/A _13409_/B VGND VGND VPWR VPWR _13409_/X sky130_fd_sc_hd__or2_4
XANTENNA__22274__B1 _24709_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14389_ _20452_/A _14382_/X _13840_/X _14384_/X VGND VGND VPWR VPWR _25138_/D sky130_fd_sc_hd__a2bb2o_4
X_17177_ _17177_/A VGND VGND VPWR VPWR _17252_/C sky130_fd_sc_hd__inv_2
XFILLER_116_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25013__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16128_ _22745_/A VGND VGND VPWR VPWR _16128_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21686__A _21686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22026__B1 _21679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16059_ _24709_/Q VGND VGND VPWR VPWR _16059_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19818_ _19817_/Y _19815_/X _19700_/X _19815_/X VGND VGND VPWR VPWR _23598_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14267__B1 _13797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19749_ _13170_/B VGND VGND VPWR VPWR _19749_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21852__C _22695_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17404__A _17404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22760_ _24751_/Q _23304_/B VGND VGND VPWR VPWR _22760_/X sky130_fd_sc_hd__or2_4
XANTENNA__18953__B1 _17424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21711_ _20592_/A _14195_/B _14463_/Y _17416_/A VGND VGND VPWR VPWR _21712_/D sky130_fd_sc_hd__o22a_4
XFILLER_38_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15767__B1 _24846_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22691_ _20877_/Y _21587_/X _16685_/Y _22442_/X VGND VGND VPWR VPWR _22691_/X sky130_fd_sc_hd__o22a_4
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24430_ _24431_/CLK _16803_/X HRESETn VGND VGND VPWR VPWR _14930_/A sky130_fd_sc_hd__dfrtp_4
X_21642_ _13780_/X VGND VGND VPWR VPWR _21816_/B sky130_fd_sc_hd__buf_2
XANTENNA__23948__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15859__A _21071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23141__A _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24361_ _24362_/CLK _17163_/X HRESETn VGND VGND VPWR VPWR _17162_/A sky130_fd_sc_hd__dfrtp_4
X_21573_ _21316_/A VGND VGND VPWR VPWR _21573_/X sky130_fd_sc_hd__buf_2
XFILLER_21_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23312_ _22534_/X _23309_/Y _23150_/X _23311_/X VGND VGND VPWR VPWR _23312_/X sky130_fd_sc_hd__a2bb2o_4
X_20524_ _24066_/Q _20519_/B _20490_/Y _20523_/X VGND VGND VPWR VPWR _20524_/X sky130_fd_sc_hd__a211o_4
XFILLER_36_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24292_ _25526_/CLK _17651_/Y HRESETn VGND VGND VPWR VPWR _24292_/Q sky130_fd_sc_hd__dfrtp_4
X_23243_ _24563_/Q _23069_/B _23005_/C VGND VGND VPWR VPWR _23243_/X sky130_fd_sc_hd__and3_4
X_20455_ _14081_/A _20455_/B VGND VGND VPWR VPWR _20455_/X sky130_fd_sc_hd__and2_4
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22804__A2 _22523_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23174_ _24427_/Q _22929_/X _22997_/X _23173_/X VGND VGND VPWR VPWR _23174_/X sky130_fd_sc_hd__a211o_4
X_20386_ _20380_/X VGND VGND VPWR VPWR _20386_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22125_ _22138_/A VGND VGND VPWR VPWR _22125_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_102_0_HCLK clkbuf_7_51_0_HCLK/X VGND VGND VPWR VPWR _24883_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__17712__A1_N _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24736__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_165_0_HCLK clkbuf_7_82_0_HCLK/X VGND VGND VPWR VPWR _23649_/CLK sky130_fd_sc_hd__clkbuf_1
X_22056_ _22055_/X _20195_/Y VGND VGND VPWR VPWR _22056_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_8_0_HCLK clkbuf_7_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21007_ _21007_/A _24841_/Q VGND VGND VPWR VPWR _21007_/X sky130_fd_sc_hd__and2_4
XANTENNA__17444__B1 _17443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13760_ _13754_/A _13758_/B _13759_/Y VGND VGND VPWR VPWR _13760_/X sky130_fd_sc_hd__o21a_4
XFILLER_90_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22958_ _22753_/X _22956_/X _22684_/X _22957_/X VGND VGND VPWR VPWR _22958_/X sky130_fd_sc_hd__o22a_4
XFILLER_56_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12711_ _12510_/Y _12713_/B _12710_/Y VGND VGND VPWR VPWR _12711_/X sky130_fd_sc_hd__o21a_4
X_21909_ _21905_/X _21908_/X _14749_/A VGND VGND VPWR VPWR _21909_/X sky130_fd_sc_hd__o21a_4
X_13691_ _13691_/A _13691_/B VGND VGND VPWR VPWR _13698_/B sky130_fd_sc_hd__or2_4
X_22889_ _23002_/A _22877_/Y _22889_/C _22889_/D VGND VGND VPWR VPWR _22889_/X sky130_fd_sc_hd__or4_4
X_12642_ _12693_/A _12642_/B VGND VGND VPWR VPWR _12645_/B sky130_fd_sc_hd__or2_4
X_15430_ _23987_/Q _14249_/A _13964_/B _15435_/A VGND VGND VPWR VPWR _15430_/X sky130_fd_sc_hd__o22a_4
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24628_ _24612_/CLK _16290_/X HRESETn VGND VGND VPWR VPWR _23247_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23296__A2 _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25524__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ _15139_/Y _15373_/A VGND VGND VPWR VPWR _15365_/B sky130_fd_sc_hd__or2_4
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ _12651_/A _24865_/Q _12651_/A _24865_/Q VGND VGND VPWR VPWR _12573_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24559_ _24557_/CLK _16477_/X HRESETn VGND VGND VPWR VPWR _16476_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18145__A _18177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17100_ _17033_/D _17091_/X VGND VGND VPWR VPWR _17100_/X sky130_fd_sc_hd__or2_4
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14312_ _14306_/X _14310_/X _25310_/Q _14311_/X VGND VGND VPWR VPWR _25164_/D sky130_fd_sc_hd__o22a_4
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15292_ _15336_/A VGND VGND VPWR VPWR _15310_/B sky130_fd_sc_hd__buf_2
X_18080_ _18080_/A _23873_/Q VGND VGND VPWR VPWR _18082_/B sky130_fd_sc_hd__or2_4
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _13914_/X VGND VGND VPWR VPWR _14244_/D sky130_fd_sc_hd__inv_2
X_17031_ _17031_/A VGND VGND VPWR VPWR _17033_/C sky130_fd_sc_hd__inv_2
XANTENNA__19121__B1 _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14174_ _14170_/Y _14173_/Y _14165_/X VGND VGND VPWR VPWR _14174_/X sky130_fd_sc_hd__o21a_4
XFILLER_98_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_61_0_HCLK clkbuf_6_30_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13125_ _24000_/Q _13124_/Y VGND VGND VPWR VPWR _13126_/B sky130_fd_sc_hd__or2_4
X_18982_ _18982_/A VGND VGND VPWR VPWR _18982_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12921__A _12936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24477__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13056_ _12988_/A _13060_/B _13055_/Y VGND VGND VPWR VPWR _25341_/D sky130_fd_sc_hd__o21a_4
X_17933_ _17955_/A _17933_/B VGND VGND VPWR VPWR _17933_/X sky130_fd_sc_hd__or2_4
X_12007_ _25299_/Q _12006_/Y _25299_/Q _12006_/Y VGND VGND VPWR VPWR _12007_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17435__B1 _16717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24406__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17864_ _17846_/X _17850_/X _17790_/A _17861_/B VGND VGND VPWR VPWR _17865_/A sky130_fd_sc_hd__a211o_4
XFILLER_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19603_ _19601_/Y _19602_/X _19553_/X _19602_/X VGND VGND VPWR VPWR _19603_/X sky130_fd_sc_hd__a2bb2o_4
X_16815_ _14971_/Y _16811_/X HWDATA[22] _16811_/X VGND VGND VPWR VPWR _24423_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17795_ _17794_/X VGND VGND VPWR VPWR _17795_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22130__A _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19534_ _22386_/A VGND VGND VPWR VPWR _19534_/Y sky130_fd_sc_hd__inv_2
X_16746_ _16745_/Y _16743_/X _15729_/X _16743_/X VGND VGND VPWR VPWR _24456_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13958_ _13958_/A _13957_/X _13958_/C _13958_/D VGND VGND VPWR VPWR _13958_/X sky130_fd_sc_hd__or4_4
XFILLER_59_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22731__A1 _22510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18935__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12909_ _12936_/A _12907_/X _12908_/X VGND VGND VPWR VPWR _12909_/X sky130_fd_sc_hd__and3_4
X_19465_ _19464_/Y _19459_/X _19420_/X _19446_/Y VGND VGND VPWR VPWR _19465_/X sky130_fd_sc_hd__a2bb2o_4
X_16677_ _22872_/A _16671_/X _16408_/X _16676_/X VGND VGND VPWR VPWR _24484_/D sky130_fd_sc_hd__a2bb2o_4
X_13889_ _24957_/Q _13920_/A _13889_/C _24954_/Q VGND VGND VPWR VPWR _13889_/X sky130_fd_sc_hd__or4_4
XFILLER_62_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18416_ _18416_/A VGND VGND VPWR VPWR _18416_/Y sky130_fd_sc_hd__inv_2
X_15628_ _15625_/Y _15626_/X _15627_/X _15626_/X VGND VGND VPWR VPWR _24885_/D sky130_fd_sc_hd__a2bb2o_4
X_19396_ _23741_/Q VGND VGND VPWR VPWR _19396_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20585__A _14394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25265__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18347_ _13190_/A _18340_/B _18344_/X VGND VGND VPWR VPWR _24190_/D sky130_fd_sc_hd__a21oi_4
X_15559_ _15559_/A VGND VGND VPWR VPWR _15559_/Y sky130_fd_sc_hd__inv_2
X_18278_ _20000_/C _18319_/B _17713_/X _18278_/D VGND VGND VPWR VPWR _18278_/X sky130_fd_sc_hd__and4_4
X_17229_ _17229_/A _17229_/B _17229_/C _17229_/D VGND VGND VPWR VPWR _17230_/D sky130_fd_sc_hd__or4_4
XANTENNA__13199__A _11964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20240_ _20240_/A VGND VGND VPWR VPWR _20240_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25127__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20171_ _22376_/B _20170_/X _20079_/X _20170_/X VGND VGND VPWR VPWR _23468_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16303__A _16288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17526__A2_N _17525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_238_0_HCLK clkbuf_8_239_0_HCLK/A VGND VGND VPWR VPWR _25330_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24147__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17426__B1 _17424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23930_ _25098_/CLK _20976_/A HRESETn VGND VGND VPWR VPWR _20977_/C sky130_fd_sc_hd__dfstp_4
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11859__A1_N _11855_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23861_ _25488_/CLK _19059_/X VGND VGND VPWR VPWR _23861_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15988__B1 _15840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19179__B1 _19133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22812_ _24551_/Q _22810_/X _22812_/C VGND VGND VPWR VPWR _22812_/X sky130_fd_sc_hd__and3_4
X_23792_ _23847_/CLK _23792_/D VGND VGND VPWR VPWR _23792_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13463__B2 _11964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18926__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25531_ _25436_/CLK _25531_/D HRESETn VGND VGND VPWR VPWR _25531_/Q sky130_fd_sc_hd__dfrtp_4
X_22743_ _21280_/B _22742_/X _21296_/X _16037_/A _21299_/X VGND VGND VPWR VPWR _22743_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_80_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12278__A _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22694__B _22298_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25462_ _23933_/CLK _12110_/X HRESETn VGND VGND VPWR VPWR _25462_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22674_ _21095_/X _22672_/X _22613_/B _22673_/X VGND VGND VPWR VPWR _22674_/X sky130_fd_sc_hd__o22a_4
X_24413_ _24413_/CLK _16835_/X HRESETn VGND VGND VPWR VPWR _24413_/Q sky130_fd_sc_hd__dfrtp_4
X_21625_ _21619_/X _21624_/X _14712_/X VGND VGND VPWR VPWR _21625_/X sky130_fd_sc_hd__o21a_4
X_25393_ _24457_/CLK _25393_/D HRESETn VGND VGND VPWR VPWR _12560_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24344_ _24330_/CLK _24344_/D HRESETn VGND VGND VPWR VPWR _24344_/Q sky130_fd_sc_hd__dfrtp_4
X_21556_ _21556_/A VGND VGND VPWR VPWR _21556_/X sky130_fd_sc_hd__buf_2
XFILLER_90_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20507_ _14205_/Y _14207_/Y _20479_/A _20479_/C VGND VGND VPWR VPWR _20507_/X sky130_fd_sc_hd__and4_4
XANTENNA__24988__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24275_ _24275_/CLK _17774_/Y HRESETn VGND VGND VPWR VPWR _24275_/Q sky130_fd_sc_hd__dfrtp_4
X_21487_ _21650_/A _19576_/Y VGND VGND VPWR VPWR _21487_/X sky130_fd_sc_hd__or2_4
XFILLER_10_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24917__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23226_ _16650_/Y _23226_/B VGND VGND VPWR VPWR _23226_/X sky130_fd_sc_hd__and2_4
X_20438_ _14063_/X _20425_/X _20429_/Y _20437_/X VGND VGND VPWR VPWR _20512_/B sky130_fd_sc_hd__a211o_4
XFILLER_10_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_48_0_HCLK clkbuf_6_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_48_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13837__A _11838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23157_ _17236_/Y _22908_/X _25381_/Q _22909_/X VGND VGND VPWR VPWR _23158_/B sky130_fd_sc_hd__a2bb2o_4
X_20369_ _21934_/B _20366_/X _19622_/A _20366_/X VGND VGND VPWR VPWR _23392_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14479__B1 _14414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22108_ _12111_/Y _21561_/X _18376_/Y _21562_/X VGND VGND VPWR VPWR _22108_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24570__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23202__A2 _22467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23088_ _22714_/X _23088_/B VGND VGND VPWR VPWR _23088_/Y sky130_fd_sc_hd__nor2_4
X_14930_ _14930_/A VGND VGND VPWR VPWR _14930_/Y sky130_fd_sc_hd__inv_2
X_22039_ _25054_/Q _19601_/Y _22036_/X _22038_/X VGND VGND VPWR VPWR _22039_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14861_ _14813_/C _14798_/X _14813_/C _14798_/X VGND VGND VPWR VPWR _14861_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15979__B1 _15758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16600_ HWDATA[9] VGND VGND VPWR VPWR _16600_/X sky130_fd_sc_hd__buf_2
X_13812_ _12095_/Y _16453_/A VGND VGND VPWR VPWR _13813_/B sky130_fd_sc_hd__or2_4
Xclkbuf_4_3_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17580_ _17580_/A _17571_/Y _17653_/B VGND VGND VPWR VPWR _17611_/B sky130_fd_sc_hd__or3_4
X_14792_ _14792_/A _13623_/A _14792_/C _14791_/X VGND VGND VPWR VPWR _14792_/X sky130_fd_sc_hd__or4_4
XFILLER_1_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22713__A1 _16130_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22885__A _22885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22713__B2 _22271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16531_ _16466_/A VGND VGND VPWR VPWR _16531_/X sky130_fd_sc_hd__buf_2
X_13743_ _13743_/A _13743_/B VGND VGND VPWR VPWR _16173_/B sky130_fd_sc_hd__or2_4
XANTENNA__17979__A _18217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19250_ _19248_/Y _19244_/X _16872_/X _19249_/X VGND VGND VPWR VPWR _23794_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16462_ _16457_/Y _16461_/X _16376_/X _16461_/X VGND VGND VPWR VPWR _16462_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13674_ _25285_/Q _13524_/X _13673_/Y VGND VGND VPWR VPWR _13674_/X sky130_fd_sc_hd__o21a_4
XFILLER_71_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15746__A3 _15745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18201_ _18201_/A _18199_/X _18200_/X VGND VGND VPWR VPWR _18201_/X sky130_fd_sc_hd__and3_4
X_15413_ _15413_/A VGND VGND VPWR VPWR _15413_/Y sky130_fd_sc_hd__inv_2
X_12625_ _25419_/Q _12625_/B VGND VGND VPWR VPWR _12625_/X sky130_fd_sc_hd__or2_4
X_19181_ _19175_/Y VGND VGND VPWR VPWR _19181_/X sky130_fd_sc_hd__buf_2
XANTENNA__15499__A _15490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16393_ HWDATA[24] VGND VGND VPWR VPWR _16393_/X sky130_fd_sc_hd__buf_2
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19342__B1 _19206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18132_ _18196_/A _18132_/B VGND VGND VPWR VPWR _18132_/X sky130_fd_sc_hd__or2_4
XANTENNA__11820__A _25517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12556_ _25406_/Q _12555_/A _12681_/A _12555_/Y VGND VGND VPWR VPWR _12557_/D sky130_fd_sc_hd__o22a_4
X_15344_ _15344_/A VGND VGND VPWR VPWR _15345_/B sky130_fd_sc_hd__inv_2
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18063_ _18196_/A _23753_/Q VGND VGND VPWR VPWR _18065_/B sky130_fd_sc_hd__or2_4
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ _12278_/B _12471_/D VGND VGND VPWR VPWR _12491_/B sky130_fd_sc_hd__or2_4
X_15275_ _15249_/A _15249_/B _15190_/A _15272_/Y VGND VGND VPWR VPWR _15276_/A sky130_fd_sc_hd__a211o_4
XFILLER_8_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15903__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17014_ _24731_/Q _17005_/Y _16066_/Y _24364_/Q VGND VGND VPWR VPWR _17014_/X sky130_fd_sc_hd__a2bb2o_4
X_14226_ _25187_/Q VGND VGND VPWR VPWR _14226_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24658__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14157_ _14129_/X _14156_/X _25123_/Q _14136_/X VGND VGND VPWR VPWR _14157_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_99_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13108_ _12993_/A _13107_/X VGND VGND VPWR VPWR _13110_/A sky130_fd_sc_hd__nand2_4
X_14088_ _13985_/B _14081_/X _14069_/X _25216_/Q _14084_/X VGND VGND VPWR VPWR _14088_/X
+ sky130_fd_sc_hd__a32o_4
X_18965_ _18965_/A VGND VGND VPWR VPWR _18965_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24240__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13039_ _12999_/D _13017_/D _12999_/B VGND VGND VPWR VPWR _13039_/X sky130_fd_sc_hd__o21a_4
X_17916_ _17915_/Y _15912_/X _17920_/C VGND VGND VPWR VPWR _17916_/X sky130_fd_sc_hd__a21o_4
XANTENNA__22401__B1 _24814_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15962__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18896_ _18894_/Y _18895_/Y _17443_/X _18895_/Y VGND VGND VPWR VPWR _18896_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17847_ _17747_/D _17792_/C VGND VGND VPWR VPWR _17848_/B sky130_fd_sc_hd__or2_4
XFILLER_93_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18620__A2 _24121_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_68_0_HCLK clkbuf_8_69_0_HCLK/A VGND VGND VPWR VPWR _23995_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17778_ _16916_/Y _17776_/A VGND VGND VPWR VPWR _17779_/C sky130_fd_sc_hd__or2_4
XANTENNA__22795__A _22795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22704__A1 _24717_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15985__A3 _15768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25446__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19517_ _22340_/B _19516_/X _11930_/X _19516_/X VGND VGND VPWR VPWR _23700_/D sky130_fd_sc_hd__a2bb2o_4
X_16729_ _16733_/A VGND VGND VPWR VPWR _16730_/A sky130_fd_sc_hd__buf_2
XANTENNA__20715__B1 _20706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17187__A2 _23072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19448_ _19444_/Y _19447_/X _19426_/X _19447_/X VGND VGND VPWR VPWR _23724_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16395__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22468__B1 _24816_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21204__A _24310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19379_ _19384_/A VGND VGND VPWR VPWR _19379_/X sky130_fd_sc_hd__buf_2
X_21410_ _21410_/A VGND VGND VPWR VPWR _23100_/A sky130_fd_sc_hd__buf_2
XFILLER_124_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22390_ _22390_/A _22390_/B VGND VGND VPWR VPWR _22390_/X sky130_fd_sc_hd__or2_4
X_21341_ _14397_/Y _14194_/A _14490_/Y _14257_/A VGND VGND VPWR VPWR _21341_/X sky130_fd_sc_hd__o22a_4
XFILLER_135_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18513__A _18460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24399__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24060_ _24496_/CLK _24060_/D HRESETn VGND VGND VPWR VPWR _24060_/Q sky130_fd_sc_hd__dfrtp_4
X_21272_ _21272_/A _21208_/X _21272_/C _21272_/D VGND VGND VPWR VPWR _21273_/A sky130_fd_sc_hd__and4_4
XFILLER_118_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20481__C _20481_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23011_ _22270_/X _23008_/X _23010_/X VGND VGND VPWR VPWR _23030_/B sky130_fd_sc_hd__and3_4
X_20223_ _20223_/A VGND VGND VPWR VPWR _20223_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21443__A1 _22792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24328__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20154_ _20161_/A VGND VGND VPWR VPWR _20154_/X sky130_fd_sc_hd__buf_2
XFILLER_104_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22689__B _22613_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20085_ _20085_/A VGND VGND VPWR VPWR _20085_/X sky130_fd_sc_hd__buf_2
XFILLER_131_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23280__A2_N _23277_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24962_ _24957_/CLK _15436_/Y HRESETn VGND VGND VPWR VPWR _13945_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_134_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22943__A1 _12849_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23913_ _24396_/CLK _23913_/D VGND VGND VPWR VPWR _18909_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_100_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14488__A _14481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24893_ _24893_/CLK _15606_/X HRESETn VGND VGND VPWR VPWR _15604_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23963__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23844_ _25316_/CLK _23844_/D VGND VGND VPWR VPWR _13180_/B sky130_fd_sc_hd__dfxtp_4
X_23775_ _23618_/CLK _19303_/X VGND VGND VPWR VPWR _13387_/B sky130_fd_sc_hd__dfxtp_4
X_20987_ _23367_/Q VGND VGND VPWR VPWR _20988_/B sky130_fd_sc_hd__inv_2
XFILLER_60_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25116__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19572__B1 _11948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25514_ _25514_/CLK _11834_/X HRESETn VGND VGND VPWR VPWR _11831_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22726_ _22726_/A _22726_/B VGND VGND VPWR VPWR _22726_/X sky130_fd_sc_hd__and2_4
XANTENNA__21114__A _21408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25445_ _25449_/CLK _12420_/X HRESETn VGND VGND VPWR VPWR _12184_/A sky130_fd_sc_hd__dfrtp_4
X_22657_ _22565_/X _22653_/Y _21045_/X _22656_/X VGND VGND VPWR VPWR _22658_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12410_ _12410_/A VGND VGND VPWR VPWR _12412_/A sky130_fd_sc_hd__buf_2
XFILLER_43_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21608_ _21608_/A _19097_/Y VGND VGND VPWR VPWR _21608_/X sky130_fd_sc_hd__or2_4
X_13390_ _13390_/A _13390_/B _13389_/X VGND VGND VPWR VPWR _13398_/B sky130_fd_sc_hd__or3_4
Xclkbuf_4_11_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_22_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_25376_ _25368_/CLK _12909_/X HRESETn VGND VGND VPWR VPWR _25376_/Q sky130_fd_sc_hd__dfrtp_4
X_22588_ _22545_/X _22587_/X _22127_/C _24853_/Q _22547_/X VGND VGND VPWR VPWR _22589_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_127_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12341_ _24824_/Q VGND VGND VPWR VPWR _12341_/Y sky130_fd_sc_hd__inv_2
X_21539_ _21275_/X _21516_/X _21522_/X _21535_/X _21538_/X VGND VGND VPWR VPWR _21539_/X
+ sky130_fd_sc_hd__o41a_4
X_24327_ _23964_/CLK _17405_/X HRESETn VGND VGND VPWR VPWR _20992_/A sky130_fd_sc_hd__dfstp_4
XFILLER_138_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12373__A2_N _24810_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15060_ _15197_/A _15194_/A VGND VGND VPWR VPWR _15070_/C sky130_fd_sc_hd__or2_4
XANTENNA__24751__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12272_ _12272_/A _12251_/X _12262_/X _12272_/D VGND VGND VPWR VPWR _12273_/B sky130_fd_sc_hd__or4_4
X_24258_ _24682_/CLK _24258_/D HRESETn VGND VGND VPWR VPWR _17752_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14670__B _13598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14011_ _13989_/X VGND VGND VPWR VPWR _14012_/C sky130_fd_sc_hd__inv_2
XANTENNA__24069__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23209_ _23190_/X _23193_/X _23197_/Y _23208_/X VGND VGND VPWR VPWR HRDATA[27] sky130_fd_sc_hd__a211o_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24189_ _24187_/CLK _24189_/D HRESETn VGND VGND VPWR VPWR _18359_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12902__C _12600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18750_ _18759_/A _18748_/X _18749_/X VGND VGND VPWR VPWR _24134_/D sky130_fd_sc_hd__and3_4
X_15962_ HWDATA[18] VGND VGND VPWR VPWR _15962_/X sky130_fd_sc_hd__buf_2
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13675__A1 _13536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_221_0_HCLK clkbuf_8_221_0_HCLK/A VGND VGND VPWR VPWR _25001_/CLK sky130_fd_sc_hd__clkbuf_1
X_17701_ _11900_/A _11871_/A _21686_/A _11899_/A VGND VGND VPWR VPWR _17702_/A sky130_fd_sc_hd__or4_4
XFILLER_49_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14913_ _14913_/A VGND VGND VPWR VPWR _14913_/Y sky130_fd_sc_hd__inv_2
X_18681_ _18681_/A VGND VGND VPWR VPWR _18682_/A sky130_fd_sc_hd__inv_2
X_15893_ _15886_/X _15887_/X _11812_/X _22623_/A _15888_/X VGND VGND VPWR VPWR _15893_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_75_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17632_ _17541_/Y _17626_/X _17601_/X _17628_/Y VGND VGND VPWR VPWR _17633_/A sky130_fd_sc_hd__a211o_4
XANTENNA__11815__A _25518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14844_ _14825_/X _14842_/Y _14802_/A _14843_/X VGND VGND VPWR VPWR _25038_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17563_ _17562_/Y _17616_/A VGND VGND VPWR VPWR _17582_/C sky130_fd_sc_hd__or2_4
X_14775_ _14764_/Y _14772_/X _14762_/C _14774_/X VGND VGND VPWR VPWR _25047_/D sky130_fd_sc_hd__o22a_4
X_11987_ _11987_/A VGND VGND VPWR VPWR _11987_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19302_ _19287_/Y VGND VGND VPWR VPWR _19302_/X sky130_fd_sc_hd__buf_2
X_16514_ _16513_/Y _16511_/X _16340_/X _16511_/X VGND VGND VPWR VPWR _16514_/X sky130_fd_sc_hd__a2bb2o_4
X_13726_ _13685_/B _13725_/Y _13721_/X _13714_/A _11656_/A VGND VGND VPWR VPWR _25272_/D
+ sky130_fd_sc_hd__a32o_4
X_17494_ _17494_/A VGND VGND VPWR VPWR _17494_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16377__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19233_ _19231_/Y _19227_/X _19232_/X _19227_/X VGND VGND VPWR VPWR _19233_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21024__A _21024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16445_ _16445_/A VGND VGND VPWR VPWR _16445_/Y sky130_fd_sc_hd__inv_2
X_13657_ _24034_/Q _13657_/B VGND VGND VPWR VPWR _13658_/B sky130_fd_sc_hd__or2_4
XFILLER_108_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16118__A _16094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12608_ _25409_/Q VGND VGND VPWR VPWR _12670_/A sky130_fd_sc_hd__inv_2
X_19164_ _18123_/B VGND VGND VPWR VPWR _19164_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16129__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24839__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16376_ HWDATA[31] VGND VGND VPWR VPWR _16376_/X sky130_fd_sc_hd__buf_2
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13588_ _13554_/X _13588_/B _13578_/X _13587_/X VGND VGND VPWR VPWR _13588_/X sky130_fd_sc_hd__or4_4
XFILLER_129_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18115_ _18080_/A _23872_/Q VGND VGND VPWR VPWR _18115_/X sky130_fd_sc_hd__or2_4
X_15327_ _15326_/X VGND VGND VPWR VPWR _24991_/D sky130_fd_sc_hd__inv_2
XANTENNA__15957__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12539_ _12539_/A VGND VGND VPWR VPWR _12539_/Y sky130_fd_sc_hd__inv_2
X_19095_ _19095_/A VGND VGND VPWR VPWR _21753_/B sky130_fd_sc_hd__inv_2
XANTENNA__22870__B1 _25373_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24492__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18046_ _18046_/A _18995_/A VGND VGND VPWR VPWR _18047_/C sky130_fd_sc_hd__or2_4
X_15258_ _15258_/A VGND VGND VPWR VPWR _15258_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24421__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14209_ _14209_/A VGND VGND VPWR VPWR _14209_/Y sky130_fd_sc_hd__inv_2
X_15189_ _15070_/X _15171_/X _15071_/A VGND VGND VPWR VPWR _15189_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21694__A _24775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_31_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16301__B1 _16300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19997_ _23533_/Q VGND VGND VPWR VPWR _19997_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18948_ _18944_/Y _18947_/X _17418_/X _18947_/X VGND VGND VPWR VPWR _23900_/D sky130_fd_sc_hd__a2bb2o_4
X_18879_ _18879_/A _18878_/X VGND VGND VPWR VPWR _18879_/X sky130_fd_sc_hd__or2_4
XFILLER_55_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20910_ _24050_/Q VGND VGND VPWR VPWR _20910_/Y sky130_fd_sc_hd__inv_2
X_21890_ _21391_/A VGND VGND VPWR VPWR _21890_/X sky130_fd_sc_hd__buf_2
XANTENNA__25280__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20841_ _13659_/B VGND VGND VPWR VPWR _20852_/B sky130_fd_sc_hd__inv_2
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18508__A _16448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19554__B1 _19553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17412__A _14807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23560_ _25264_/CLK _19921_/X VGND VGND VPWR VPWR _23560_/Q sky130_fd_sc_hd__dfxtp_4
X_20772_ _13120_/A _13120_/B _20772_/C _13120_/D VGND VGND VPWR VPWR _20772_/X sky130_fd_sc_hd__or4_4
XFILLER_35_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22511_ _22508_/X _22511_/B VGND VGND VPWR VPWR _22511_/Y sky130_fd_sc_hd__nor2_4
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23491_ _23434_/CLK _20109_/X VGND VGND VPWR VPWR _23491_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12929__B1 _12874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22442_ _23069_/B VGND VGND VPWR VPWR _22442_/X sky130_fd_sc_hd__buf_2
XFILLER_91_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25230_ _24955_/CLK _25230_/D HRESETn VGND VGND VPWR VPWR scl_oen_o_S5 sky130_fd_sc_hd__dfstp_4
XANTENNA__13197__A3 _13195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21113__B1 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17868__B1 _16955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24509__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25161_ _25305_/CLK _25161_/D HRESETn VGND VGND VPWR VPWR _25161_/Q sky130_fd_sc_hd__dfrtp_4
X_22373_ _22369_/X _22372_/X _14677_/X VGND VGND VPWR VPWR _22373_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__22861__B1 _16029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_113_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_227_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24112_ _24136_/CLK _18867_/Y HRESETn VGND VGND VPWR VPWR pwm_S7 sky130_fd_sc_hd__dfrtp_4
X_21324_ _21293_/A VGND VGND VPWR VPWR _22592_/B sky130_fd_sc_hd__buf_2
X_25092_ _25093_/CLK _25092_/D HRESETn VGND VGND VPWR VPWR _21709_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16540__B1 _16366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24043_ _24496_/CLK _20881_/X HRESETn VGND VGND VPWR VPWR _20879_/A sky130_fd_sc_hd__dfrtp_4
X_21255_ _21252_/A _20144_/Y VGND VGND VPWR VPWR _21255_/X sky130_fd_sc_hd__or2_4
XFILLER_135_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12291__A _12291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20206_ _20205_/Y _20203_/X _19797_/A _20203_/X VGND VGND VPWR VPWR _23454_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21186_ _21186_/A _21186_/B _21186_/C VGND VGND VPWR VPWR _21186_/X sky130_fd_sc_hd__and3_4
XFILLER_132_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20137_ _23480_/Q VGND VGND VPWR VPWR _21772_/B sky130_fd_sc_hd__inv_2
XFILLER_131_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25368__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20068_ _20064_/X _18326_/X _11838_/A _23507_/Q _20066_/X VGND VGND VPWR VPWR _20068_/X
+ sky130_fd_sc_hd__a32o_4
X_24945_ _24945_/CLK _24945_/D HRESETn VGND VGND VPWR VPWR _24945_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_86_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11910_ _11871_/A _11700_/X _11902_/X _11909_/Y VGND VGND VPWR VPWR _11910_/X sky130_fd_sc_hd__a211o_4
XFILLER_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12890_ _12749_/A _12890_/B VGND VGND VPWR VPWR _12890_/X sky130_fd_sc_hd__or2_4
XFILLER_73_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24876_ _23805_/CLK _15689_/Y HRESETn VGND VGND VPWR VPWR _24876_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_51_0_HCLK clkbuf_8_51_0_HCLK/A VGND VGND VPWR VPWR _25081_/CLK sky130_fd_sc_hd__clkbuf_1
X_11841_ HWDATA[5] VGND VGND VPWR VPWR _11842_/A sky130_fd_sc_hd__buf_2
X_23827_ _23884_/CLK _23827_/D VGND VGND VPWR VPWR _19157_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_26_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19545__B1 _19407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17322__A _17254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13850__A _23990_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11772_ _11770_/Y _11768_/X _11771_/X _11768_/X VGND VGND VPWR VPWR _25530_/D sky130_fd_sc_hd__a2bb2o_4
X_14560_ _14560_/A _14560_/B VGND VGND VPWR VPWR _14560_/X sky130_fd_sc_hd__or2_4
XFILLER_14_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23758_ _23869_/CLK _19350_/X VGND VGND VPWR VPWR _19348_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_92_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13511_ _25296_/Q VGND VGND VPWR VPWR _13511_/Y sky130_fd_sc_hd__inv_2
X_22709_ _24856_/Q _22707_/X _21103_/A _22708_/X VGND VGND VPWR VPWR _22710_/C sky130_fd_sc_hd__a211o_4
X_14491_ _14490_/Y _14488_/X _14470_/X _14488_/X VGND VGND VPWR VPWR _25102_/D sky130_fd_sc_hd__a2bb2o_4
X_23689_ _23689_/CLK _23689_/D VGND VGND VPWR VPWR _23689_/Q sky130_fd_sc_hd__dfxtp_4
X_16230_ _16230_/A VGND VGND VPWR VPWR _16230_/Y sky130_fd_sc_hd__inv_2
X_13442_ _13156_/X _13440_/X _13441_/X VGND VGND VPWR VPWR _13442_/X sky130_fd_sc_hd__and3_4
XANTENNA__24932__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25428_ _25425_/CLK _25428_/D HRESETn VGND VGND VPWR VPWR _12202_/A sky130_fd_sc_hd__dfrtp_4
X_13373_ _13373_/A _13373_/B VGND VGND VPWR VPWR _13374_/C sky130_fd_sc_hd__or2_4
X_16161_ _21513_/A VGND VGND VPWR VPWR _16161_/Y sky130_fd_sc_hd__inv_2
X_25359_ _25330_/CLK _25359_/D HRESETn VGND VGND VPWR VPWR _25359_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_5_24_0_HCLK_A clkbuf_4_12_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15112_ _24576_/Q VGND VGND VPWR VPWR _15112_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12324_ _24814_/Q VGND VGND VPWR VPWR _12324_/Y sky130_fd_sc_hd__inv_2
X_16092_ _16092_/A VGND VGND VPWR VPWR _16092_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12255_ _23210_/A VGND VGND VPWR VPWR _12255_/Y sky130_fd_sc_hd__inv_2
X_15043_ _25019_/Q _15042_/Y _25019_/Q _15042_/Y VGND VGND VPWR VPWR _15047_/B sky130_fd_sc_hd__a2bb2o_4
X_19920_ _23560_/Q VGND VGND VPWR VPWR _19920_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19851_ _19851_/A VGND VGND VPWR VPWR _19851_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12186_ _12178_/X _12186_/B _12183_/X _12185_/X VGND VGND VPWR VPWR _12186_/X sky130_fd_sc_hd__or4_4
Xclkbuf_5_18_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_122_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24581__CLK _24581_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18802_ _18786_/C _18786_/D VGND VGND VPWR VPWR _18803_/B sky130_fd_sc_hd__or2_4
X_19782_ _23610_/Q VGND VGND VPWR VPWR _19782_/Y sky130_fd_sc_hd__inv_2
X_16994_ _16994_/A VGND VGND VPWR VPWR _17130_/A sky130_fd_sc_hd__inv_2
XANTENNA__16401__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18733_ _18733_/A VGND VGND VPWR VPWR _18733_/X sky130_fd_sc_hd__buf_2
XFILLER_49_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12250__A2_N _24750_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15945_ _15938_/X VGND VGND VPWR VPWR _15945_/X sky130_fd_sc_hd__buf_2
XANTENNA__21019__A _21019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25038__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18664_ _24530_/Q _18705_/B _16613_/Y _24117_/Q VGND VGND VPWR VPWR _18666_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15876_ _12772_/Y _15872_/X _11767_/X _15872_/X VGND VGND VPWR VPWR _15876_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16598__B1 _16340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21591__B1 _21587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17615_ _17562_/Y _17617_/B _17614_/Y VGND VGND VPWR VPWR _17615_/X sky130_fd_sc_hd__o21a_4
XFILLER_92_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14827_ _25042_/Q _14804_/A _14819_/C _14806_/B VGND VGND VPWR VPWR _14827_/X sky130_fd_sc_hd__o22a_4
X_18595_ _18475_/D _18496_/X _18498_/X _18592_/Y VGND VGND VPWR VPWR _18595_/X sky130_fd_sc_hd__a211o_4
XANTENNA__18856__A1_N _24558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12265__A2_N _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17546_ _11850_/Y _17573_/A _11860_/A _17578_/C VGND VGND VPWR VPWR _17550_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12084__B1 _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14758_ _21622_/A VGND VGND VPWR VPWR _21608_/A sky130_fd_sc_hd__buf_2
X_13709_ _13698_/B _13707_/X _13708_/Y _13703_/X _25279_/Q VGND VGND VPWR VPWR _13709_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_36_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17477_ _17477_/A VGND VGND VPWR VPWR _17477_/Y sky130_fd_sc_hd__inv_2
X_14689_ _14689_/A VGND VGND VPWR VPWR _14752_/A sky130_fd_sc_hd__buf_2
X_19216_ _18222_/B VGND VGND VPWR VPWR _19216_/Y sky130_fd_sc_hd__inv_2
X_16428_ _15086_/Y _16426_/X _16340_/X _16426_/X VGND VGND VPWR VPWR _24577_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24673__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19147_ _19146_/Y _19144_/X _19056_/X _19144_/X VGND VGND VPWR VPWR _19147_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21646__A1 _21634_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24602__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16359_ _16359_/A VGND VGND VPWR VPWR _16359_/X sky130_fd_sc_hd__buf_2
XFILLER_9_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19078_ _19075_/Y _19076_/X _19077_/X _19076_/X VGND VGND VPWR VPWR _19078_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16522__B1 _16521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18029_ _18066_/A _19317_/A VGND VGND VPWR VPWR _18031_/B sky130_fd_sc_hd__or2_4
XFILLER_99_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21040_ _21040_/A _21026_/X _21040_/C VGND VGND VPWR VPWR _21040_/X sky130_fd_sc_hd__and3_4
XFILLER_99_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24070__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13639__A1 _14620_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16311__A _16288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25461__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23020__B1 _22090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22991_ _22088_/A VGND VGND VPWR VPWR _23133_/A sky130_fd_sc_hd__buf_2
X_24730_ _24712_/CLK _16008_/X HRESETn VGND VGND VPWR VPWR _24730_/Q sky130_fd_sc_hd__dfrtp_4
X_21942_ _21942_/A _19523_/Y VGND VGND VPWR VPWR _21942_/X sky130_fd_sc_hd__or2_4
XANTENNA__16589__B1 _16231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_38_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_77_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21873_ _12819_/X _21872_/X _17745_/A _21422_/X VGND VGND VPWR VPWR _21873_/X sky130_fd_sc_hd__a2bb2o_4
X_24661_ _24162_/CLK _16198_/X HRESETn VGND VGND VPWR VPWR _23200_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _20816_/X VGND VGND VPWR VPWR _20824_/X sky130_fd_sc_hd__buf_2
XANTENNA__17142__A _17038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23612_ _23609_/CLK _23612_/D VGND VGND VPWR VPWR _23612_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12075__B1 _11833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21590__A2_N _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24592_ _24995_/CLK _16392_/X HRESETn VGND VGND VPWR VPWR _24592_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20755_ _13119_/A _20750_/X _20754_/X VGND VGND VPWR VPWR _20755_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23543_ _24309_/CLK _19965_/X VGND VGND VPWR VPWR _19963_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_50_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12286__A _12199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23087__B1 _12321_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23474_ _23562_/CLK _23474_/D VGND VGND VPWR VPWR _20153_/A sky130_fd_sc_hd__dfxtp_4
X_20686_ _20678_/X VGND VGND VPWR VPWR _20686_/X sky130_fd_sc_hd__buf_2
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_HCLK clkbuf_3_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22425_ _22425_/A VGND VGND VPWR VPWR _22425_/X sky130_fd_sc_hd__buf_2
XANTENNA__24343__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25213_ _24322_/CLK _25213_/D HRESETn VGND VGND VPWR VPWR _14003_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_104_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22356_ _14682_/B _19773_/Y VGND VGND VPWR VPWR _22356_/X sky130_fd_sc_hd__or2_4
X_25144_ _25141_/CLK _25144_/D HRESETn VGND VGND VPWR VPWR _25144_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21307_ _24030_/Q _21302_/X _21305_/X _21306_/X VGND VGND VPWR VPWR _21307_/X sky130_fd_sc_hd__a211o_4
X_25075_ _25081_/CLK _14603_/X HRESETn VGND VGND VPWR VPWR _13559_/A sky130_fd_sc_hd__dfrtp_4
X_22287_ _22287_/A _22286_/X VGND VGND VPWR VPWR _22287_/X sky130_fd_sc_hd__and2_4
XFILLER_136_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12040_ _12040_/A VGND VGND VPWR VPWR _12040_/Y sky130_fd_sc_hd__inv_2
X_24026_ _24026_/CLK _20806_/X HRESETn VGND VGND VPWR VPWR _20804_/A sky130_fd_sc_hd__dfrtp_4
X_21238_ _14691_/A VGND VGND VPWR VPWR _21238_/X sky130_fd_sc_hd__buf_2
XANTENNA__18266__B1 _16852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17317__A _17254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21169_ _21173_/A _19997_/Y VGND VGND VPWR VPWR _21169_/X sky130_fd_sc_hd__or2_4
XANTENNA__23038__B _23037_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16221__A _22809_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13991_ _13999_/A _25227_/Q _13990_/X VGND VGND VPWR VPWR _14040_/C sky130_fd_sc_hd__or3_4
XFILLER_59_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15730_ _15728_/X _15713_/X _15729_/X _24865_/Q _15711_/X VGND VGND VPWR VPWR _15730_/X
+ sky130_fd_sc_hd__a32o_4
X_12942_ _12819_/X _12941_/X VGND VGND VPWR VPWR _12959_/B sky130_fd_sc_hd__or2_4
XFILLER_20_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21781__B _21504_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24928_ _24926_/CLK _15507_/X HRESETn VGND VGND VPWR VPWR _15506_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15661_ _12095_/A _16453_/A VGND VGND VPWR VPWR _15662_/D sky130_fd_sc_hd__or2_4
X_12873_ _12881_/A _12873_/B _12873_/C VGND VGND VPWR VPWR _12873_/X sky130_fd_sc_hd__and3_4
X_24859_ _24847_/CLK _15738_/X HRESETn VGND VGND VPWR VPWR _12559_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_65_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17400_ _17402_/B VGND VGND VPWR VPWR _17401_/A sky130_fd_sc_hd__inv_2
X_14612_ _25070_/Q _14599_/X _13770_/X _14560_/B VGND VGND VPWR VPWR _25070_/D sky130_fd_sc_hd__o22a_4
X_11824_ _11824_/A VGND VGND VPWR VPWR _11824_/Y sky130_fd_sc_hd__inv_2
X_18380_ _18379_/Y _18377_/X _18381_/A _18377_/X VGND VGND VPWR VPWR _18380_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14999__A2_N _16785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15592_ _24898_/Q VGND VGND VPWR VPWR _15592_/Y sky130_fd_sc_hd__inv_2
XPHY_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17250_/A _17331_/B VGND VGND VPWR VPWR _17331_/X sky130_fd_sc_hd__or2_4
XFILLER_60_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14543_ _14006_/X _14043_/Y _14543_/C VGND VGND VPWR VPWR _14547_/C sky130_fd_sc_hd__or3_4
XANTENNA__17987__A _17995_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11753_/Y _11751_/X _11754_/X _11751_/X VGND VGND VPWR VPWR _25535_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12196__A _21065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _17262_/A VGND VGND VPWR VPWR _17263_/B sky130_fd_sc_hd__inv_2
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14474_ _14474_/A VGND VGND VPWR VPWR _14474_/Y sky130_fd_sc_hd__inv_2
X_11686_ _24221_/Q VGND VGND VPWR VPWR _11686_/Y sky130_fd_sc_hd__inv_2
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19001_ _19000_/Y _18998_/X _18955_/X _18998_/X VGND VGND VPWR VPWR _23881_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16213_ _16211_/Y _16212_/X _15955_/X _16212_/X VGND VGND VPWR VPWR _16213_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24084__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13425_ _13457_/A _13425_/B _13424_/X VGND VGND VPWR VPWR _13429_/B sky130_fd_sc_hd__and3_4
X_17193_ _22899_/A _17192_/A _16315_/Y _17254_/C VGND VGND VPWR VPWR _17193_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15300__A _24973_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24013__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16144_ _16125_/X VGND VGND VPWR VPWR _16144_/X sky130_fd_sc_hd__buf_2
X_13356_ _13452_/A _13356_/B VGND VGND VPWR VPWR _13357_/C sky130_fd_sc_hd__or2_4
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12307_ _12992_/A _12305_/Y _12306_/Y _24833_/Q VGND VGND VPWR VPWR _12313_/B sky130_fd_sc_hd__a2bb2o_4
X_16075_ _16075_/A VGND VGND VPWR VPWR _16075_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13287_ _13227_/A VGND VGND VPWR VPWR _13392_/A sky130_fd_sc_hd__buf_2
X_15026_ _15219_/B _24450_/Q _14903_/X _15025_/Y VGND VGND VPWR VPWR _15033_/B sky130_fd_sc_hd__a2bb2o_4
X_19903_ _21669_/B _19902_/X _19629_/X _19902_/X VGND VGND VPWR VPWR _19903_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18257__B1 _16717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12238_ _12238_/A VGND VGND VPWR VPWR _12238_/X sky130_fd_sc_hd__buf_2
XFILLER_64_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23250__B1 _16916_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12169_ _12123_/Y _12168_/Y SCLK_S3 _12167_/X VGND VGND VPWR VPWR _12169_/X sky130_fd_sc_hd__o22a_4
X_19834_ _21745_/B _19829_/X _19790_/X _19829_/X VGND VGND VPWR VPWR _19834_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16977_ _24727_/Q _24384_/Q _16014_/Y _16976_/Y VGND VGND VPWR VPWR _16977_/X sky130_fd_sc_hd__o22a_4
X_19765_ _23615_/Q VGND VGND VPWR VPWR _19765_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25292__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22787__B _22873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15928_ _15674_/X _15925_/B VGND VGND VPWR VPWR _15928_/X sky130_fd_sc_hd__or2_4
X_18716_ _18715_/X VGND VGND VPWR VPWR _18716_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21691__B _22998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19696_ _19696_/A VGND VGND VPWR VPWR _19696_/Y sky130_fd_sc_hd__inv_2
X_18647_ _24136_/Q VGND VGND VPWR VPWR _18647_/X sky130_fd_sc_hd__buf_2
X_15859_ _21071_/A VGND VGND VPWR VPWR _23035_/A sky130_fd_sc_hd__buf_2
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23305__A1 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23305__B2 _21067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24854__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18578_ _18521_/A VGND VGND VPWR VPWR _18582_/C sky130_fd_sc_hd__buf_2
XFILLER_101_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17529_ _11860_/A _17578_/C _25512_/Q _17528_/Y VGND VGND VPWR VPWR _17529_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20540_ _14446_/Y _20533_/X _14452_/X _20539_/X VGND VGND VPWR VPWR _20541_/A sky130_fd_sc_hd__a211o_4
XFILLER_71_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15806__A1_N _12321_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21212__A _21015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20471_ _20468_/Y _20469_/X _20517_/A VGND VGND VPWR VPWR _24072_/D sky130_fd_sc_hd__a21o_4
XANTENNA__16306__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22210_ _14693_/A _22208_/X _22209_/X VGND VGND VPWR VPWR _22210_/X sky130_fd_sc_hd__and3_4
XFILLER_118_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22292__A1 _23281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23190_ _23114_/A _23190_/B _23183_/X _23189_/X VGND VGND VPWR VPWR _23190_/X sky130_fd_sc_hd__or4_4
XFILLER_106_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22141_ _22141_/A _21085_/A VGND VGND VPWR VPWR _22141_/X sky130_fd_sc_hd__or2_4
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15849__A2 _15713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22072_ _21618_/A _20084_/Y VGND VGND VPWR VPWR _22072_/X sky130_fd_sc_hd__or2_4
XANTENNA__20055__B1 _19790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21023_ _21826_/A VGND VGND VPWR VPWR _21024_/A sky130_fd_sc_hd__buf_2
XANTENNA__19996__B1 _19995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16274__A2 _15993_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20070__A3 _15836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14285__A1 _23428_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19385__A2_N _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22974_ _22973_/X VGND VGND VPWR VPWR _22974_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24713_ _24318_/CLK _24713_/D HRESETn VGND VGND VPWR VPWR _24713_/Q sky130_fd_sc_hd__dfrtp_4
X_21925_ _22009_/A VGND VGND VPWR VPWR _21945_/A sky130_fd_sc_hd__buf_2
XANTENNA__24595__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24644_ _24643_/CLK _24644_/D HRESETn VGND VGND VPWR VPWR _22539_/A sky130_fd_sc_hd__dfrtp_4
X_21856_ _15671_/A VGND VGND VPWR VPWR _23082_/B sky130_fd_sc_hd__buf_2
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24524__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _13137_/C VGND VGND VPWR VPWR _20807_/Y sky130_fd_sc_hd__inv_2
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21787_ _21649_/A _21785_/X _21786_/X VGND VGND VPWR VPWR _21787_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_125_0_HCLK clkbuf_7_62_0_HCLK/X VGND VGND VPWR VPWR _24977_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24575_ _24572_/CLK _16431_/X HRESETn VGND VGND VPWR VPWR _24575_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_188_0_HCLK clkbuf_7_94_0_HCLK/X VGND VGND VPWR VPWR _25526_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23526_ _23550_/CLK _23526_/D VGND VGND VPWR VPWR _23526_/Q sky130_fd_sc_hd__dfxtp_4
X_20738_ _20740_/A VGND VGND VPWR VPWR _20738_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15537__B2 _15535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20669_ _20663_/A _20666_/Y _20667_/Y _14281_/X _20668_/X VGND VGND VPWR VPWR _20669_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23457_ _23609_/CLK _20199_/X VGND VGND VPWR VPWR _20198_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12744__A _12859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ _13225_/A VGND VGND VPWR VPWR _13379_/A sky130_fd_sc_hd__buf_2
X_22408_ _22278_/X _22406_/X _22280_/X _22407_/X VGND VGND VPWR VPWR _22409_/B sky130_fd_sc_hd__o22a_4
X_14190_ _16371_/A _14190_/B VGND VGND VPWR VPWR _14195_/A sky130_fd_sc_hd__or2_4
X_23388_ _23388_/CLK _23388_/D VGND VGND VPWR VPWR _20377_/A sky130_fd_sc_hd__dfxtp_4
X_13141_ _24839_/Q VGND VGND VPWR VPWR _13141_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15037__A2_N _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25127_ _25101_/CLK _14427_/X HRESETn VGND VGND VPWR VPWR _25127_/Q sky130_fd_sc_hd__dfstp_4
X_22339_ _21929_/A _22339_/B VGND VGND VPWR VPWR _22341_/B sky130_fd_sc_hd__or2_4
XFILLER_109_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25383__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13072_ _12347_/Y _13071_/X VGND VGND VPWR VPWR _13073_/A sky130_fd_sc_hd__or2_4
XFILLER_112_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25058_ _25044_/CLK _14673_/X HRESETn VGND VGND VPWR VPWR _25058_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20046__B1 _19777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12023_ _12023_/A VGND VGND VPWR VPWR _12023_/Y sky130_fd_sc_hd__inv_2
X_16900_ _16900_/A VGND VGND VPWR VPWR _16900_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25312__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24009_ _24041_/CLK _20733_/X HRESETn VGND VGND VPWR VPWR _13132_/A sky130_fd_sc_hd__dfrtp_4
X_17880_ _17748_/Y _17878_/X _17879_/Y VGND VGND VPWR VPWR _17880_/X sky130_fd_sc_hd__o21a_4
XFILLER_120_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16831_ _16829_/Y _16825_/X _15745_/X _16830_/X VGND VGND VPWR VPWR _16831_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23157__A1_N _17236_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19550_ _19549_/Y _19544_/X _19389_/X _19544_/X VGND VGND VPWR VPWR _23688_/D sky130_fd_sc_hd__a2bb2o_4
X_16762_ _16761_/Y _16759_/X _15743_/X _16759_/X VGND VGND VPWR VPWR _16762_/X sky130_fd_sc_hd__a2bb2o_4
X_13974_ _14042_/A VGND VGND VPWR VPWR _13975_/A sky130_fd_sc_hd__inv_2
X_18501_ _18503_/B VGND VGND VPWR VPWR _18506_/B sky130_fd_sc_hd__inv_2
XANTENNA__22400__B _22266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15713_ _15713_/A VGND VGND VPWR VPWR _15713_/X sky130_fd_sc_hd__buf_2
X_12925_ _12927_/B VGND VGND VPWR VPWR _12926_/B sky130_fd_sc_hd__inv_2
X_19481_ _21807_/B _19476_/X _11948_/X _19476_/X VGND VGND VPWR VPWR _19481_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17214__B2 _17252_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16693_ _22598_/A _16688_/X _15752_/X _16688_/X VGND VGND VPWR VPWR _24477_/D sky130_fd_sc_hd__a2bb2o_4
X_18432_ _16234_/Y _18467_/A _16234_/Y _18467_/A VGND VGND VPWR VPWR _18432_/X sky130_fd_sc_hd__a2bb2o_4
X_15644_ _15526_/Y _11731_/C _11731_/D _14433_/A VGND VGND VPWR VPWR _15648_/A sky130_fd_sc_hd__or4_4
XFILLER_33_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_21_0_HCLK clkbuf_7_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12856_ _12602_/A _12855_/X VGND VGND VPWR VPWR _12856_/X sky130_fd_sc_hd__or2_4
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24265__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_84_0_HCLK clkbuf_7_85_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_84_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11807_ _25520_/Q VGND VGND VPWR VPWR _11807_/Y sky130_fd_sc_hd__inv_2
X_18363_ _18363_/A _18353_/Y VGND VGND VPWR VPWR _18363_/Y sky130_fd_sc_hd__nor2_4
X_15575_ _15563_/A VGND VGND VPWR VPWR _15575_/X sky130_fd_sc_hd__buf_2
X_12787_ _25357_/Q VGND VGND VPWR VPWR _12845_/B sky130_fd_sc_hd__inv_2
XPHY_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _17306_/X _17312_/X _17313_/X VGND VGND VPWR VPWR _24349_/D sky130_fd_sc_hd__and3_4
X_14526_ _21709_/A _14510_/X _21542_/A _14505_/X VGND VGND VPWR VPWR _14526_/X sky130_fd_sc_hd__o22a_4
XPHY_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _21066_/A VGND VGND VPWR VPWR _22913_/A sky130_fd_sc_hd__buf_2
X_18294_ _18291_/X _18301_/B VGND VGND VPWR VPWR _18295_/A sky130_fd_sc_hd__and2_4
XANTENNA__22128__A _15625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16536__A1_N _16535_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17245_ _17244_/Y _17199_/Y _17245_/C VGND VGND VPWR VPWR _17245_/X sky130_fd_sc_hd__or3_4
X_14457_ _14456_/Y _14454_/X _14414_/X _14454_/X VGND VGND VPWR VPWR _14457_/X sky130_fd_sc_hd__a2bb2o_4
X_11669_ _11669_/A VGND VGND VPWR VPWR _11669_/Y sky130_fd_sc_hd__inv_2
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _13440_/A _23372_/Q VGND VGND VPWR VPWR _13410_/B sky130_fd_sc_hd__or2_4
XFILLER_122_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22274__A1 _22271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17176_ _24609_/Q _17350_/C _16295_/Y _17236_/A VGND VGND VPWR VPWR _17176_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22274__B2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14388_ _25138_/Q VGND VGND VPWR VPWR _20452_/A sky130_fd_sc_hd__inv_2
XFILLER_122_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16127_ _16124_/Y _16126_/X _11796_/X _16126_/X VGND VGND VPWR VPWR _16127_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12762__B2 _24772_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13339_ _13260_/X _13337_/X _13338_/X VGND VGND VPWR VPWR _13339_/X sky130_fd_sc_hd__and3_4
XANTENNA__22981__A1_N _12285_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21686__B _21816_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16058_ _16056_/Y _16052_/X _16057_/X _16052_/X VGND VGND VPWR VPWR _16058_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20037__B1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25053__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15009_ _14915_/A _24441_/Q _15251_/B _15008_/Y VGND VGND VPWR VPWR _15012_/C sky130_fd_sc_hd__o22a_4
XFILLER_97_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18245__A3 _16600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22798__A _22798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19817_ _19817_/A VGND VGND VPWR VPWR _19817_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19748_ _19747_/Y _19743_/X _19658_/X _19729_/Y VGND VGND VPWR VPWR _23621_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21537__B1 _25357_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19679_ _19678_/Y _19676_/X _19462_/X _19676_/X VGND VGND VPWR VPWR _19679_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20111__A _20105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11733__A _11733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21710_ _14423_/Y _14223_/A _14446_/Y _15462_/A VGND VGND VPWR VPWR _21710_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15767__A1 _15749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22690_ _22505_/X _22688_/X _21950_/A _22689_/Y VGND VGND VPWR VPWR _22690_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16964__B1 _16033_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20760__B2 _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21641_ _22531_/B _21640_/X _13565_/Y _22531_/B VGND VGND VPWR VPWR _21641_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18516__A _24168_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21572_ _14937_/Y _21570_/X _21316_/A _21571_/X VGND VGND VPWR VPWR _21572_/X sky130_fd_sc_hd__o22a_4
X_24360_ _24362_/CLK _17165_/Y HRESETn VGND VGND VPWR VPWR _17043_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20523_ _20468_/Y _20522_/X _24073_/Q VGND VGND VPWR VPWR _20523_/X sky130_fd_sc_hd__o21a_4
XFILLER_138_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23311_ _22545_/X _23310_/X _22127_/C _11706_/A _22547_/X VGND VGND VPWR VPWR _23311_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_18_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24291_ _24305_/CLK _17658_/X HRESETn VGND VGND VPWR VPWR _24291_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23988__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20454_ _20443_/A _20439_/X _20454_/C VGND VGND VPWR VPWR _20455_/B sky130_fd_sc_hd__and3_4
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22319__A1_N _14807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23242_ _23242_/A _22884_/B VGND VGND VPWR VPWR _23245_/B sky130_fd_sc_hd__or2_4
XFILLER_105_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23917__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23173_ _24459_/Q _22998_/X _23172_/X VGND VGND VPWR VPWR _23173_/X sky130_fd_sc_hd__o21a_4
X_20385_ _23385_/Q VGND VGND VPWR VPWR _20385_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22124_ _24471_/Q _22836_/B VGND VGND VPWR VPWR _22124_/X sky130_fd_sc_hd__or2_4
X_22055_ _21253_/A VGND VGND VPWR VPWR _22055_/X sky130_fd_sc_hd__buf_2
XFILLER_121_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21006_ _21006_/A _21006_/B VGND VGND VPWR VPWR _21006_/X sky130_fd_sc_hd__and2_4
XFILLER_43_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24776__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21117__A _24919_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24705__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22957_ _16115_/Y _22513_/B _15931_/B _11780_/Y _22846_/X VGND VGND VPWR VPWR _22957_/X
+ sky130_fd_sc_hd__o32a_4
X_12710_ _12510_/Y _12713_/B _12653_/X VGND VGND VPWR VPWR _12710_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_43_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21908_ _21890_/X _21906_/X _21907_/X VGND VGND VPWR VPWR _21908_/X sky130_fd_sc_hd__and3_4
X_13690_ _13690_/A _13689_/X VGND VGND VPWR VPWR _13691_/B sky130_fd_sc_hd__or2_4
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22888_ _23065_/A _22884_/X _22888_/C VGND VGND VPWR VPWR _22889_/D sky130_fd_sc_hd__and3_4
X_12641_ _12641_/A VGND VGND VPWR VPWR _12641_/Y sky130_fd_sc_hd__inv_2
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24627_ _24612_/CLK _16292_/X HRESETn VGND VGND VPWR VPWR _24627_/Q sky130_fd_sc_hd__dfrtp_4
X_21839_ _16451_/A _21836_/X _21839_/C VGND VGND VPWR VPWR _21862_/A sky130_fd_sc_hd__and3_4
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15360_ _15130_/Y _15352_/B VGND VGND VPWR VPWR _15373_/A sky130_fd_sc_hd__or2_4
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _12659_/A VGND VGND VPWR VPWR _12651_/A sky130_fd_sc_hd__inv_2
XANTENNA__12441__B1 _12394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24558_ _24557_/CLK _16480_/X HRESETn VGND VGND VPWR VPWR _24558_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ _13644_/X VGND VGND VPWR VPWR _14311_/X sky130_fd_sc_hd__buf_2
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23509_ _25055_/CLK _20062_/X VGND VGND VPWR VPWR _20061_/A sky130_fd_sc_hd__dfxtp_4
X_15291_ _15387_/B VGND VGND VPWR VPWR _15336_/A sky130_fd_sc_hd__buf_2
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24489_ _24447_/CLK _24489_/D HRESETn VGND VGND VPWR VPWR _24489_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17030_ _17030_/A VGND VGND VPWR VPWR _17105_/A sky130_fd_sc_hd__inv_2
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14242_ _14241_/Y _14236_/X _13810_/X _14224_/A VGND VGND VPWR VPWR _14242_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15785__A _15931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14173_ _14173_/A _14173_/B VGND VGND VPWR VPWR _14173_/Y sky130_fd_sc_hd__nor2_4
X_13124_ _13123_/X VGND VGND VPWR VPWR _13124_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23205__B1 _23172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18981_ _18980_/Y _18978_/X _18961_/X _18978_/X VGND VGND VPWR VPWR _18981_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11818__A _11818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13055_ _12988_/A _13060_/B _13031_/X VGND VGND VPWR VPWR _13055_/Y sky130_fd_sc_hd__a21oi_4
X_17932_ _17929_/A VGND VGND VPWR VPWR _17955_/A sky130_fd_sc_hd__buf_2
XFILLER_79_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19830__A2_N _19824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12006_ _12006_/A VGND VGND VPWR VPWR _12006_/Y sky130_fd_sc_hd__inv_2
X_17863_ _17874_/A _17863_/B _17863_/C VGND VGND VPWR VPWR _17863_/X sky130_fd_sc_hd__and3_4
XANTENNA__18632__B1 _16599_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19602_ _19587_/X VGND VGND VPWR VPWR _19602_/X sky130_fd_sc_hd__buf_2
X_16814_ _16813_/Y _16811_/X _15729_/X _16811_/X VGND VGND VPWR VPWR _24424_/D sky130_fd_sc_hd__a2bb2o_4
X_17794_ _16909_/Y _17794_/B VGND VGND VPWR VPWR _17794_/X sky130_fd_sc_hd__or2_4
XANTENNA__23226__B _23226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16745_ _16745_/A VGND VGND VPWR VPWR _16745_/Y sky130_fd_sc_hd__inv_2
X_19533_ _21174_/B _19528_/X _19488_/X _19528_/A VGND VGND VPWR VPWR _19533_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24446__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13957_ _13945_/A _13957_/B VGND VGND VPWR VPWR _13957_/X sky130_fd_sc_hd__or2_4
XANTENNA__22731__A2 _22728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21534__A3 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12908_ _12849_/C _12905_/X VGND VGND VPWR VPWR _12908_/X sky130_fd_sc_hd__or2_4
X_19464_ _18206_/B VGND VGND VPWR VPWR _19464_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16676_ _16664_/A VGND VGND VPWR VPWR _16676_/X sky130_fd_sc_hd__buf_2
X_13888_ _13945_/A VGND VGND VPWR VPWR _13953_/A sky130_fd_sc_hd__buf_2
X_15627_ _16528_/A VGND VGND VPWR VPWR _15627_/X sky130_fd_sc_hd__buf_2
X_18415_ _23242_/A _18414_/A _16191_/Y _18481_/B VGND VGND VPWR VPWR _18422_/A sky130_fd_sc_hd__o22a_4
XANTENNA__23242__A _23242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12839_ _12979_/A VGND VGND VPWR VPWR _12881_/A sky130_fd_sc_hd__buf_2
X_19395_ _19394_/Y _19392_/X _19349_/X _19392_/X VGND VGND VPWR VPWR _23742_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12174__A1_N SSn_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18346_ _13191_/A _18344_/X _18345_/Y VGND VGND VPWR VPWR _24191_/D sky130_fd_sc_hd__o21a_4
X_15558_ _15548_/X _15552_/Y _15553_/X _23318_/A _15560_/A VGND VGND VPWR VPWR _15558_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_128_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14509_ _20441_/A _14507_/X _14502_/X _14508_/Y VGND VGND VPWR VPWR _25098_/D sky130_fd_sc_hd__a211o_4
X_18277_ _24205_/Q VGND VGND VPWR VPWR _18278_/D sky130_fd_sc_hd__buf_2
Xclkbuf_8_171_0_HCLK clkbuf_7_85_0_HCLK/X VGND VGND VPWR VPWR _24926_/CLK sky130_fd_sc_hd__clkbuf_1
X_15489_ _24064_/D VGND VGND VPWR VPWR _15516_/A sky130_fd_sc_hd__inv_2
X_17228_ _16349_/Y _17168_/A _16358_/Y _24331_/Q VGND VGND VPWR VPWR _17229_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21697__A _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_28_0_HCLK clkbuf_8_29_0_HCLK/A VGND VGND VPWR VPWR _23933_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__14724__A2 _14675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12189__A1_N _12440_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23049__A1_N _17257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25234__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17159_ _16985_/Y _17159_/B VGND VGND VPWR VPWR _17160_/B sky130_fd_sc_hd__nand2_4
X_20170_ _20182_/A VGND VGND VPWR VPWR _20170_/X sky130_fd_sc_hd__buf_2
XFILLER_115_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20106__A _20105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23860_ _25316_/CLK _19064_/X VGND VGND VPWR VPWR _23860_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12757__A1_N _12843_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24187__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22811_ _15854_/X VGND VGND VPWR VPWR _22812_/C sky130_fd_sc_hd__buf_2
X_23791_ _23846_/CLK _19257_/X VGND VGND VPWR VPWR _19255_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24116__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25530_ _24759_/CLK _25530_/D HRESETn VGND VGND VPWR VPWR _25530_/Q sky130_fd_sc_hd__dfrtp_4
X_22742_ _24614_/Q _22592_/B VGND VGND VPWR VPWR _22742_/X sky130_fd_sc_hd__or2_4
XANTENNA__12278__B _12278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25461_ _25461_/CLK _12112_/X HRESETn VGND VGND VPWR VPWR _25461_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22673_ _11697_/Y _21950_/A _13569_/Y _22505_/A VGND VGND VPWR VPWR _22673_/X sky130_fd_sc_hd__o22a_4
XFILLER_40_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24412_ _24998_/CLK _24412_/D HRESETn VGND VGND VPWR VPWR _24412_/Q sky130_fd_sc_hd__dfrtp_4
X_21624_ _21624_/A _21621_/X _21624_/C VGND VGND VPWR VPWR _21624_/X sky130_fd_sc_hd__and3_4
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22486__B2 _22915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25392_ _24457_/CLK _25392_/D HRESETn VGND VGND VPWR VPWR _25392_/Q sky130_fd_sc_hd__dfrtp_4
X_24343_ _24345_/CLK _24343_/D HRESETn VGND VGND VPWR VPWR _17250_/A sky130_fd_sc_hd__dfrtp_4
X_21555_ _21548_/Y _21549_/Y _21552_/Y _21554_/Y VGND VGND VPWR VPWR _21555_/X sky130_fd_sc_hd__or4_4
X_20506_ _20506_/A _14282_/X _14281_/X VGND VGND VPWR VPWR _20506_/X sky130_fd_sc_hd__and3_4
X_21486_ _21455_/A VGND VGND VPWR VPWR _21650_/A sky130_fd_sc_hd__buf_2
X_24274_ _24267_/CLK _24274_/D HRESETn VGND VGND VPWR VPWR _16916_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_119_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20437_ _20451_/A _20458_/A _20437_/C _20436_/X VGND VGND VPWR VPWR _20437_/X sky130_fd_sc_hd__or4_4
XANTENNA__19077__A _16442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23225_ _23223_/X _23224_/X _22132_/A VGND VGND VPWR VPWR _23225_/X sky130_fd_sc_hd__or3_4
XFILLER_10_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20368_ _20368_/A VGND VGND VPWR VPWR _21934_/B sky130_fd_sc_hd__inv_2
X_23156_ _12290_/A _22980_/X _17740_/A _22906_/X VGND VGND VPWR VPWR _23156_/X sky130_fd_sc_hd__a2bb2o_4
X_22107_ _13505_/Y _12097_/X _12033_/Y _21562_/X VGND VGND VPWR VPWR _22107_/X sky130_fd_sc_hd__o22a_4
XFILLER_122_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24957__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23087_ _12207_/Y _22426_/X _22712_/X _12321_/Y _22840_/X VGND VGND VPWR VPWR _23088_/B
+ sky130_fd_sc_hd__o32a_4
X_20299_ _20298_/Y VGND VGND VPWR VPWR _20299_/X sky130_fd_sc_hd__buf_2
X_22038_ _22038_/A _19606_/Y _22037_/X VGND VGND VPWR VPWR _22038_/X sky130_fd_sc_hd__and3_4
XFILLER_130_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14860_ _14845_/X _14859_/Y _15467_/A _14811_/X VGND VGND VPWR VPWR _14860_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13811_ _13808_/Y _13804_/X _13810_/X _13804_/X VGND VGND VPWR VPWR _25258_/D sky130_fd_sc_hd__a2bb2o_4
X_14791_ _14663_/D _14790_/X _14663_/D _14790_/X VGND VGND VPWR VPWR _14791_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23989_ _23989_/CLK _20672_/X HRESETn VGND VGND VPWR VPWR _23989_/Q sky130_fd_sc_hd__dfrtp_4
X_16530_ _21837_/A VGND VGND VPWR VPWR _16530_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22713__A2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13742_ _13742_/A VGND VGND VPWR VPWR _13743_/B sky130_fd_sc_hd__inv_2
XFILLER_1_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20686__A _20678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16461_ _16461_/A VGND VGND VPWR VPWR _16461_/X sky130_fd_sc_hd__buf_2
XFILLER_16_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13673_ _13673_/A VGND VGND VPWR VPWR _13673_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18200_ _18168_/A _23445_/Q VGND VGND VPWR VPWR _18200_/X sky130_fd_sc_hd__or2_4
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15412_ _15389_/A _15388_/X _15409_/Y _15339_/X VGND VGND VPWR VPWR _15413_/A sky130_fd_sc_hd__a211o_4
X_12624_ _12626_/B VGND VGND VPWR VPWR _12625_/B sky130_fd_sc_hd__inv_2
X_19180_ _19180_/A VGND VGND VPWR VPWR _19180_/Y sky130_fd_sc_hd__inv_2
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16392_ _16391_/Y _16389_/X _16300_/X _16389_/X VGND VGND VPWR VPWR _16392_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18131_ _17963_/X _18130_/X _24232_/Q _18021_/X VGND VGND VPWR VPWR _24232_/D sky130_fd_sc_hd__o22a_4
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15343_ _15346_/A _15338_/X _15343_/C VGND VGND VPWR VPWR _15343_/X sky130_fd_sc_hd__and3_4
XFILLER_8_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17995__A _17995_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ _12555_/A VGND VGND VPWR VPWR _12555_/Y sky130_fd_sc_hd__inv_2
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_244_0_HCLK clkbuf_8_245_0_HCLK/A VGND VGND VPWR VPWR _24431_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18062_ _13610_/A VGND VGND VPWR VPWR _18196_/A sky130_fd_sc_hd__buf_2
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15274_ _15282_/A _15267_/B _15273_/X VGND VGND VPWR VPWR _15274_/X sky130_fd_sc_hd__and3_4
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12486_ _12485_/X VGND VGND VPWR VPWR _25428_/D sky130_fd_sc_hd__inv_2
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17013_ _15999_/Y _17022_/A _15999_/Y _17022_/A VGND VGND VPWR VPWR _17013_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14225_ _14218_/Y _14224_/X _13835_/X _14224_/X VGND VGND VPWR VPWR _25188_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12932__A _12799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14156_ _14100_/A _14100_/B _14100_/A _14100_/B VGND VGND VPWR VPWR _14156_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18853__B1 _16508_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13107_ _13107_/A _13106_/X VGND VGND VPWR VPWR _13107_/X sky130_fd_sc_hd__or2_4
XANTENNA__19715__A _15766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24698__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14087_ _25216_/Q _14081_/X _14078_/X _13983_/X _14084_/X VGND VGND VPWR VPWR _14087_/X
+ sky130_fd_sc_hd__a32o_4
X_18964_ _18963_/Y _18960_/X _18940_/X _18960_/X VGND VGND VPWR VPWR _23894_/D sky130_fd_sc_hd__a2bb2o_4
X_13038_ _13038_/A _13038_/B _13037_/X VGND VGND VPWR VPWR _25345_/D sky130_fd_sc_hd__and3_4
X_17915_ _13541_/X VGND VGND VPWR VPWR _17915_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22401__A1 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24627__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18895_ _18895_/A _21116_/A VGND VGND VPWR VPWR _18895_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22141__A _22141_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17846_ _17846_/A VGND VGND VPWR VPWR _17846_/X sky130_fd_sc_hd__buf_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24280__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14989_ _14961_/X _24448_/Q _14961_/X _24448_/Q VGND VGND VPWR VPWR _14996_/B sky130_fd_sc_hd__a2bb2o_4
X_17777_ _16916_/A _17776_/Y VGND VGND VPWR VPWR _17779_/B sky130_fd_sc_hd__or2_4
XFILLER_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22704__A2 _22407_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19516_ _19528_/A VGND VGND VPWR VPWR _19516_/X sky130_fd_sc_hd__buf_2
XFILLER_47_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16728_ _16728_/A _16728_/B VGND VGND VPWR VPWR _16733_/A sky130_fd_sc_hd__nor2_4
X_16659_ _23120_/A _16658_/X _16300_/X _16658_/X VGND VGND VPWR VPWR _24491_/D sky130_fd_sc_hd__a2bb2o_4
X_19447_ _19446_/Y VGND VGND VPWR VPWR _19447_/X sky130_fd_sc_hd__buf_2
XFILLER_35_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25486__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22468__A1 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_54_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19378_ _19377_/X VGND VGND VPWR VPWR _19384_/A sky130_fd_sc_hd__buf_2
XANTENNA__22468__B2 _22467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25415__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18329_ _19728_/A _17462_/Y _19683_/C VGND VGND VPWR VPWR _18329_/X sky130_fd_sc_hd__or3_4
X_21340_ _21339_/X VGND VGND VPWR VPWR _21340_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21220__A _21220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21271_ _21261_/X _21268_/X _21270_/X VGND VGND VPWR VPWR _21272_/D sky130_fd_sc_hd__a21o_4
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17726__A1_N _17722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12842__A _12842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20222_ _20221_/Y _20217_/X _19740_/X _20217_/X VGND VGND VPWR VPWR _23448_/D sky130_fd_sc_hd__a2bb2o_4
X_23010_ _24725_/Q _21021_/X _21050_/X _23009_/X VGND VGND VPWR VPWR _23010_/X sky130_fd_sc_hd__a211o_4
XFILLER_104_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22640__A1 _12799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20153_ _20153_/A VGND VGND VPWR VPWR _22075_/B sky130_fd_sc_hd__inv_2
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23147__A _16295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24368__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20084_ _23498_/Q VGND VGND VPWR VPWR _20084_/Y sky130_fd_sc_hd__inv_2
X_24961_ _24957_/CLK _15439_/X HRESETn VGND VGND VPWR VPWR _24961_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22051__A _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14769__A _13588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20403__B1 _19755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23912_ _23847_/CLK _18912_/X VGND VGND VPWR VPWR _23912_/Q sky130_fd_sc_hd__dfxtp_4
X_24892_ _24893_/CLK _15608_/X HRESETn VGND VGND VPWR VPWR _24892_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16997__A1_N _16039_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23843_ _23441_/CLK _19110_/X VGND VGND VPWR VPWR _13206_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12289__A _12244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15830__B1 _15758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19021__B1 _18993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23774_ _23618_/CLK _19305_/X VGND VGND VPWR VPWR _13419_/B sky130_fd_sc_hd__dfxtp_4
X_20986_ _14214_/Y _14196_/X VGND VGND VPWR VPWR _23959_/D sky130_fd_sc_hd__and2_4
XFILLER_53_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25513_ _25514_/CLK _11839_/X HRESETn VGND VGND VPWR VPWR _25513_/Q sky130_fd_sc_hd__dfrtp_4
X_22725_ _22574_/A _22722_/X _22725_/C VGND VGND VPWR VPWR _22725_/X sky130_fd_sc_hd__and3_4
XFILLER_41_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25444_ _25449_/CLK _12422_/Y HRESETn VGND VGND VPWR VPWR _12206_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23932__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22656_ _15709_/A _22655_/X _22130_/C _25520_/Q _22677_/B VGND VGND VPWR VPWR _22656_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21607_ _21629_/A _21607_/B VGND VGND VPWR VPWR _21607_/X sky130_fd_sc_hd__or2_4
XANTENNA__21131__A1 _25475_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25375_ _25368_/CLK _12911_/Y HRESETn VGND VGND VPWR VPWR _25375_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22587_ _24783_/Q _22587_/B VGND VGND VPWR VPWR _22587_/X sky130_fd_sc_hd__or2_4
XFILLER_51_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21131__B2 _12059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14149__B1 _25126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12340_ _12301_/X _12313_/X _12340_/C _12339_/X VGND VGND VPWR VPWR _12382_/A sky130_fd_sc_hd__or4_4
X_24326_ _23964_/CLK _17406_/X HRESETn VGND VGND VPWR VPWR _24326_/Q sky130_fd_sc_hd__dfstp_4
X_21538_ _21536_/X _21538_/B _21095_/X VGND VGND VPWR VPWR _21538_/X sky130_fd_sc_hd__or3_4
XFILLER_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12271_ _12271_/A _12271_/B _12271_/C _12271_/D VGND VGND VPWR VPWR _12272_/D sky130_fd_sc_hd__or4_4
Xclkbuf_8_11_0_HCLK clkbuf_7_5_0_HCLK/X VGND VGND VPWR VPWR _23562_/CLK sky130_fd_sc_hd__clkbuf_1
X_24257_ _24682_/CLK _17844_/Y HRESETn VGND VGND VPWR VPWR _24257_/Q sky130_fd_sc_hd__dfrtp_4
X_21469_ _21469_/A _21461_/X _21468_/X VGND VGND VPWR VPWR _21469_/X sky130_fd_sc_hd__or3_4
XFILLER_88_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14010_ _14006_/A _13999_/X _14010_/C VGND VGND VPWR VPWR _14010_/X sky130_fd_sc_hd__or3_4
Xclkbuf_8_74_0_HCLK clkbuf_8_75_0_HCLK/A VGND VGND VPWR VPWR _25101_/CLK sky130_fd_sc_hd__clkbuf_1
X_23208_ _23208_/A _23199_/Y _23203_/X _23208_/D VGND VGND VPWR VPWR _23208_/X sky130_fd_sc_hd__or4_4
X_24188_ _24187_/CLK _24188_/D HRESETn VGND VGND VPWR VPWR _24188_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19535__A _13595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24791__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23139_ _23114_/X _23117_/X _23124_/Y _23138_/X VGND VGND VPWR VPWR HRDATA[25] sky130_fd_sc_hd__a211o_4
XFILLER_68_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15961_ _12214_/Y _15954_/X _15959_/X _15960_/X VGND VGND VPWR VPWR _15961_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24720__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14912_ _15067_/A VGND VGND VPWR VPWR _15219_/A sky130_fd_sc_hd__buf_2
X_17700_ _13771_/X _11709_/B _17700_/C _17447_/X VGND VGND VPWR VPWR _17700_/X sky130_fd_sc_hd__or4_4
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24038__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15892_ _15886_/X _15887_/X _11809_/A _22651_/A _15888_/X VGND VGND VPWR VPWR _24785_/D
+ sky130_fd_sc_hd__a32o_4
X_18680_ _18680_/A _18680_/B _18678_/Y _18680_/D VGND VGND VPWR VPWR _18680_/X sky130_fd_sc_hd__or4_4
XANTENNA__16074__B1 _15840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14843_ _14824_/X VGND VGND VPWR VPWR _14843_/X sky130_fd_sc_hd__buf_2
X_17631_ _17642_/A _17629_/X _17631_/C VGND VGND VPWR VPWR _24299_/D sky130_fd_sc_hd__and3_4
XFILLER_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15821__B1 _24821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17562_ _17562_/A VGND VGND VPWR VPWR _17562_/Y sky130_fd_sc_hd__inv_2
X_14774_ _25046_/Q _25045_/Q _14776_/B VGND VGND VPWR VPWR _14774_/X sky130_fd_sc_hd__and3_4
XFILLER_112_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11986_ _11654_/A _11987_/A _11978_/Y _11985_/Y VGND VGND VPWR VPWR _11986_/X sky130_fd_sc_hd__o22a_4
X_16513_ _24544_/Q VGND VGND VPWR VPWR _16513_/Y sky130_fd_sc_hd__inv_2
X_19301_ _13387_/B VGND VGND VPWR VPWR _19301_/Y sky130_fd_sc_hd__inv_2
X_13725_ _11656_/Y _13684_/B VGND VGND VPWR VPWR _13725_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__19563__B2 _19562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17493_ _11706_/Y _24309_/Q _11706_/Y _24309_/Q VGND VGND VPWR VPWR _17497_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21370__A1 _14620_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12927__A _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11843__A1_N _11840_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11831__A _11831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16444_ _15125_/Y _16375_/A _16266_/X _16375_/A VGND VGND VPWR VPWR _16444_/X sky130_fd_sc_hd__a2bb2o_4
X_19232_ _16786_/X VGND VGND VPWR VPWR _19232_/X sky130_fd_sc_hd__buf_2
X_13656_ _13656_/A _13656_/B VGND VGND VPWR VPWR _13657_/B sky130_fd_sc_hd__or2_4
XFILLER_90_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12607_ _12517_/Y _12656_/A VGND VGND VPWR VPWR _12620_/C sky130_fd_sc_hd__or2_4
X_19163_ _19162_/Y _19160_/X _19071_/X _19160_/X VGND VGND VPWR VPWR _23825_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18441__A1_N _16199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16375_ _16375_/A VGND VGND VPWR VPWR _16375_/X sky130_fd_sc_hd__buf_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13587_ _13581_/X _13583_/X _13585_/X _13587_/D VGND VGND VPWR VPWR _13587_/X sky130_fd_sc_hd__or4_4
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18114_ _17928_/X _18114_/B _18113_/X VGND VGND VPWR VPWR _18114_/X sky130_fd_sc_hd__and3_4
X_15326_ _15309_/A _15325_/X _15318_/A _15322_/B VGND VGND VPWR VPWR _15326_/X sky130_fd_sc_hd__a211o_4
X_12538_ _25412_/Q VGND VGND VPWR VPWR _12656_/A sky130_fd_sc_hd__inv_2
X_19094_ _21888_/B _19091_/X _16876_/X _19091_/X VGND VGND VPWR VPWR _23849_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22870__B2 _22288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22136__A _21525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18045_ _18221_/A _18045_/B VGND VGND VPWR VPWR _18045_/X sky130_fd_sc_hd__or2_4
XFILLER_117_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15257_ _15251_/C _15256_/X _15190_/A _15253_/B VGND VGND VPWR VPWR _15258_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24879__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12469_ _12281_/X _12509_/B VGND VGND VPWR VPWR _12469_/X sky130_fd_sc_hd__or2_4
XANTENNA__12662__A _12631_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14208_ _14207_/Y _14199_/X _13797_/X _14201_/X VGND VGND VPWR VPWR _14208_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18826__B1 _24539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24808__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15188_ _15198_/A _15186_/X _15188_/C VGND VGND VPWR VPWR _15188_/X sky130_fd_sc_hd__and3_4
XFILLER_98_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14139_ _14117_/A _14117_/B _14117_/A _14117_/B VGND VGND VPWR VPWR _14139_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21694__B _22998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19996_ _21479_/B _19991_/X _19995_/X _19991_/X VGND VGND VPWR VPWR _19996_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24461__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18947_ _18946_/Y VGND VGND VPWR VPWR _18947_/X sky130_fd_sc_hd__buf_2
XFILLER_67_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18878_ _20574_/A _20571_/A VGND VGND VPWR VPWR _18878_/X sky130_fd_sc_hd__or2_4
XFILLER_66_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16065__B1 _16064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17829_ _17829_/A VGND VGND VPWR VPWR _24261_/D sky130_fd_sc_hd__inv_2
XFILLER_94_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19003__B1 _18977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20840_ _20839_/X VGND VGND VPWR VPWR _20840_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16080__A3 _15927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20771_ _13120_/A VGND VGND VPWR VPWR _20771_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22510_ _22510_/A VGND VGND VPWR VPWR _22511_/B sky130_fd_sc_hd__buf_2
XFILLER_50_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23490_ _23609_/CLK _20112_/X VGND VGND VPWR VPWR _20110_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22441_ _22441_/A VGND VGND VPWR VPWR _22441_/X sky130_fd_sc_hd__buf_2
XANTENNA__22310__B1 _25427_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25160_ _25305_/CLK _25160_/D HRESETn VGND VGND VPWR VPWR _25160_/Q sky130_fd_sc_hd__dfrtp_4
X_22372_ _21763_/A _22370_/X _22371_/X VGND VGND VPWR VPWR _22372_/X sky130_fd_sc_hd__and3_4
XANTENNA__22861__B2 _22480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24111_ _25199_/CLK _24111_/D HRESETn VGND VGND VPWR VPWR _20974_/A sky130_fd_sc_hd__dfstp_4
X_21323_ _21323_/A VGND VGND VPWR VPWR _21323_/X sky130_fd_sc_hd__buf_2
X_25091_ _25137_/CLK _25091_/D HRESETn VGND VGND VPWR VPWR _21542_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16540__B2 _16461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21254_ _21250_/A _21254_/B _21254_/C VGND VGND VPWR VPWR _21254_/X sky130_fd_sc_hd__and3_4
XFILLER_102_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24549__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24042_ _24496_/CLK _20876_/X HRESETn VGND VGND VPWR VPWR _13663_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20205_ _20205_/A VGND VGND VPWR VPWR _20205_/Y sky130_fd_sc_hd__inv_2
X_21185_ _21185_/A _20040_/Y VGND VGND VPWR VPWR _21186_/C sky130_fd_sc_hd__or2_4
XANTENNA__19355__A _19354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20136_ _21906_/B _20133_/X _20089_/X _20133_/X VGND VGND VPWR VPWR _20136_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24131__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20067_ _20064_/X _18326_/X _13835_/A _23508_/Q _20066_/X VGND VGND VPWR VPWR _20067_/X
+ sky130_fd_sc_hd__a32o_4
X_24944_ _24943_/CLK _24944_/D HRESETn VGND VGND VPWR VPWR _24944_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_86_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24875_ _23805_/CLK _15697_/X HRESETn VGND VGND VPWR VPWR _15680_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15803__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11840_ _25512_/Q VGND VGND VPWR VPWR _11840_/Y sky130_fd_sc_hd__inv_2
X_23826_ _23826_/CLK _23826_/D VGND VGND VPWR VPWR _19159_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23341__A2 _21979_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25337__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11771_ HWDATA[23] VGND VGND VPWR VPWR _11771_/X sky130_fd_sc_hd__buf_2
XFILLER_60_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23757_ _23722_/CLK _19352_/X VGND VGND VPWR VPWR _18214_/B sky130_fd_sc_hd__dfxtp_4
X_20969_ _20969_/A VGND VGND VPWR VPWR _20970_/B sky130_fd_sc_hd__inv_2
XANTENNA__12747__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13510_ _13509_/Y _13507_/X _11853_/X _13507_/X VGND VGND VPWR VPWR _13510_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22708_ _22708_/A _21859_/B _21859_/C VGND VGND VPWR VPWR _22708_/X sky130_fd_sc_hd__and3_4
X_14490_ _25102_/Q VGND VGND VPWR VPWR _14490_/Y sky130_fd_sc_hd__inv_2
X_23688_ _23689_/CLK _23688_/D VGND VGND VPWR VPWR _23688_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13441_ _13345_/A _18965_/A VGND VGND VPWR VPWR _13441_/X sky130_fd_sc_hd__or2_4
X_25427_ _25385_/CLK _12490_/X HRESETn VGND VGND VPWR VPWR _25427_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22639_ _17753_/Y _22821_/A _12235_/X _22429_/A VGND VGND VPWR VPWR _22639_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16160_ _16159_/Y _16157_/X _15474_/X _16157_/X VGND VGND VPWR VPWR _16160_/X sky130_fd_sc_hd__a2bb2o_4
X_13372_ _13303_/A _13372_/B VGND VGND VPWR VPWR _13372_/X sky130_fd_sc_hd__or2_4
XFILLER_10_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25358_ _25356_/CLK _25358_/D HRESETn VGND VGND VPWR VPWR _25358_/Q sky130_fd_sc_hd__dfrtp_4
X_15111_ _15111_/A VGND VGND VPWR VPWR _15299_/A sky130_fd_sc_hd__inv_2
X_12323_ _25329_/Q VGND VGND VPWR VPWR _13096_/A sky130_fd_sc_hd__inv_2
X_24309_ _24309_/CLK _17588_/X HRESETn VGND VGND VPWR VPWR _24309_/Q sky130_fd_sc_hd__dfrtp_4
X_16091_ _16090_/Y _16088_/X _11746_/X _16088_/X VGND VGND VPWR VPWR _16091_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24972__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25289_ _25054_/CLK _25289_/D HRESETn VGND VGND VPWR VPWR _25289_/Q sky130_fd_sc_hd__dfstp_4
X_15042_ _24457_/Q VGND VGND VPWR VPWR _15042_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12254_ _25424_/Q VGND VGND VPWR VPWR _12278_/C sky130_fd_sc_hd__inv_2
XANTENNA__22604__A1 _12842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24901__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19850_ _19849_/Y _19847_/X _19780_/X _19847_/X VGND VGND VPWR VPWR _23587_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19265__A _19264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12185_ _12277_/A _24760_/Q _12277_/A _24760_/Q VGND VGND VPWR VPWR _12185_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19481__B1 _11948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18801_ _18800_/X VGND VGND VPWR VPWR _18801_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19781_ _22215_/B _19776_/X _19780_/X _19776_/X VGND VGND VPWR VPWR _19781_/X sky130_fd_sc_hd__a2bb2o_4
X_16993_ _17162_/A VGND VGND VPWR VPWR _16993_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18732_ _18738_/A _18730_/X _18731_/X VGND VGND VPWR VPWR _24138_/D sky130_fd_sc_hd__and3_4
XFILLER_95_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19233__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15944_ HWDATA[27] VGND VGND VPWR VPWR _15944_/X sky130_fd_sc_hd__buf_2
XFILLER_77_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15875_ _15850_/X _15857_/X _15725_/X _24797_/Q _15864_/X VGND VGND VPWR VPWR _15875_/X
+ sky130_fd_sc_hd__a32o_4
X_18663_ _18654_/Y VGND VGND VPWR VPWR _18705_/B sky130_fd_sc_hd__buf_2
XANTENNA__21591__A1 _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14826_ _14809_/A VGND VGND VPWR VPWR _14831_/A sky130_fd_sc_hd__buf_2
X_17614_ _17562_/Y _17617_/B _17590_/X VGND VGND VPWR VPWR _17614_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18594_ _18585_/X _18594_/B _18582_/C VGND VGND VPWR VPWR _18594_/X sky130_fd_sc_hd__and3_4
XFILLER_52_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25078__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11782__A1_N _11780_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14757_ _21385_/A VGND VGND VPWR VPWR _21622_/A sky130_fd_sc_hd__buf_2
X_17545_ _17538_/X _17540_/X _17545_/C _17545_/D VGND VGND VPWR VPWR _17551_/C sky130_fd_sc_hd__or4_4
X_11969_ _11967_/D VGND VGND VPWR VPWR _11969_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25007__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13708_ _13691_/A _13691_/B VGND VGND VPWR VPWR _13708_/Y sky130_fd_sc_hd__nand2_4
X_17476_ _17476_/A _17449_/X VGND VGND VPWR VPWR _17477_/A sky130_fd_sc_hd__or2_4
X_14688_ _21245_/A VGND VGND VPWR VPWR _14689_/A sky130_fd_sc_hd__buf_2
X_19215_ _19214_/Y _19211_/X _19191_/X _19211_/X VGND VGND VPWR VPWR _23806_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13639_ _14620_/D _13633_/X _13638_/X VGND VGND VPWR VPWR _25289_/D sky130_fd_sc_hd__a21oi_4
X_16427_ _16425_/Y _16426_/X _16242_/X _16426_/X VGND VGND VPWR VPWR _16427_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16358_ _24602_/Q VGND VGND VPWR VPWR _16358_/Y sky130_fd_sc_hd__inv_2
X_19146_ _23830_/Q VGND VGND VPWR VPWR _19146_/Y sky130_fd_sc_hd__inv_2
X_15309_ _15309_/A _15331_/A _15309_/C _15308_/X VGND VGND VPWR VPWR _15309_/X sky130_fd_sc_hd__or4_4
XFILLER_118_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20854__B1 _20845_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16289_ _16288_/X VGND VGND VPWR VPWR _16289_/X sky130_fd_sc_hd__buf_2
X_19077_ _16442_/A VGND VGND VPWR VPWR _19077_/X sky130_fd_sc_hd__buf_2
XANTENNA__12392__A _12385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18028_ _17996_/A VGND VGND VPWR VPWR _18066_/A sky130_fd_sc_hd__buf_2
XANTENNA__14533__B1 _25101_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24642__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16286__B1 _16285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19979_ _22238_/B _19974_/X _19978_/X _19974_/X VGND VGND VPWR VPWR _23539_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15208__A _15246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22990_ _23056_/A _22990_/B VGND VGND VPWR VPWR _22990_/Y sky130_fd_sc_hd__nor2_4
XFILLER_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16038__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21941_ _17717_/A _21941_/B VGND VGND VPWR VPWR _21941_/X sky130_fd_sc_hd__or2_4
XFILLER_27_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24660_ _24654_/CLK _16201_/X HRESETn VGND VGND VPWR VPWR _23165_/A sky130_fd_sc_hd__dfrtp_4
X_21872_ _21009_/X VGND VGND VPWR VPWR _21872_/X sky130_fd_sc_hd__buf_2
XFILLER_83_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25430__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _23434_/CLK _19781_/X VGND VGND VPWR VPWR _23611_/Q sky130_fd_sc_hd__dfxtp_4
X_20823_ _20823_/A VGND VGND VPWR VPWR _20823_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24591_ _24995_/CLK _24591_/D HRESETn VGND VGND VPWR VPWR _24591_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17538__B1 _25517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16039__A _24717_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23542_ _23550_/CLK _19967_/X VGND VGND VPWR VPWR _23542_/Q sky130_fd_sc_hd__dfxtp_4
X_20754_ _20749_/Y _20745_/Y _20754_/C VGND VGND VPWR VPWR _20754_/X sky130_fd_sc_hd__and3_4
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16210__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12286__B _12286_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23087__A1 _12207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23473_ _23496_/CLK _20157_/X VGND VGND VPWR VPWR _23473_/Q sky130_fd_sc_hd__dfxtp_4
X_20685_ _20685_/A VGND VGND VPWR VPWR _20685_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18254__A _18254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_24_0_HCLK clkbuf_4_12_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_49_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25212_ _25093_/CLK _14121_/X HRESETn VGND VGND VPWR VPWR _25212_/Q sky130_fd_sc_hd__dfrtp_4
X_22424_ _22424_/A _22423_/X VGND VGND VPWR VPWR _22424_/Y sky130_fd_sc_hd__nor2_4
XFILLER_104_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25143_ _25141_/CLK _25143_/D HRESETn VGND VGND VPWR VPWR _25143_/Q sky130_fd_sc_hd__dfrtp_4
X_22355_ _21890_/X _22353_/X _22354_/X VGND VGND VPWR VPWR _22355_/X sky130_fd_sc_hd__and3_4
XFILLER_100_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21306_ _21306_/A VGND VGND VPWR VPWR _21306_/X sky130_fd_sc_hd__buf_2
XANTENNA__24383__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25074_ _25246_/CLK _25074_/D HRESETn VGND VGND VPWR VPWR _13582_/A sky130_fd_sc_hd__dfrtp_4
X_22286_ _21413_/X _22284_/X _22396_/C _12514_/A _22540_/A VGND VGND VPWR VPWR _22286_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_105_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19085__A _19084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24312__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24025_ _24025_/CLK _24025_/D HRESETn VGND VGND VPWR VPWR _20799_/A sky130_fd_sc_hd__dfrtp_4
X_21237_ _21250_/A _21235_/X _21236_/X VGND VGND VPWR VPWR _21237_/X sky130_fd_sc_hd__and3_4
XANTENNA__19463__B1 _19462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12550__A2 _24851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21168_ _21184_/A _21168_/B VGND VGND VPWR VPWR _21170_/B sky130_fd_sc_hd__or2_4
XANTENNA__20024__A _20036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_148_0_HCLK clkbuf_7_74_0_HCLK/X VGND VGND VPWR VPWR _24252_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_59_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20119_ _20117_/Y _20118_/X _20096_/X _20118_/X VGND VGND VPWR VPWR _20119_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19215__B1 _19191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13990_ _13997_/A _13990_/B _13990_/C _25221_/Q VGND VGND VPWR VPWR _13990_/X sky130_fd_sc_hd__or4_4
X_21099_ _17242_/A _21095_/X _21098_/X VGND VGND VPWR VPWR _21099_/X sky130_fd_sc_hd__o21a_4
XFILLER_63_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25518__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12941_ _12941_/A _12979_/B VGND VGND VPWR VPWR _12941_/X sky130_fd_sc_hd__or2_4
X_24927_ _24930_/CLK _15509_/X HRESETn VGND VGND VPWR VPWR _11729_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_73_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15660_ _15643_/Y _15655_/X _15647_/X _20812_/A _15659_/X VGND VGND VPWR VPWR _24878_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_65_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12872_ _12864_/A _12869_/X VGND VGND VPWR VPWR _12873_/C sky130_fd_sc_hd__or2_4
XFILLER_46_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24858_ _24865_/CLK _24858_/D HRESETn VGND VGND VPWR VPWR _24858_/Q sky130_fd_sc_hd__dfrtp_4
X_14611_ _14560_/X _14610_/X _14557_/X _14602_/X _14610_/A VGND VGND VPWR VPWR _14611_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11823_ _11820_/Y _11816_/X _11822_/X _11816_/X VGND VGND VPWR VPWR _11823_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23809_ _23805_/CLK _23809_/D VGND VGND VPWR VPWR _18094_/B sky130_fd_sc_hd__dfxtp_4
X_15591_ _15590_/Y _15588_/X _11784_/X _15588_/X VGND VGND VPWR VPWR _24899_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12477__A _12220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17529__B1 _25512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24789_ _24785_/CLK _24789_/D HRESETn VGND VGND VPWR VPWR _12792_/A sky130_fd_sc_hd__dfrtp_4
X_17330_ _17330_/A VGND VGND VPWR VPWR _17331_/B sky130_fd_sc_hd__inv_2
XANTENNA__19568__A2_N _19562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25100__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14535_/Y _14073_/B _20459_/B VGND VGND VPWR VPWR _14542_/X sky130_fd_sc_hd__o21a_4
XFILLER_18_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ HWDATA[28] VGND VGND VPWR VPWR _11754_/X sky130_fd_sc_hd__buf_2
XFILLER_60_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16201__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17194_/Y _17261_/B _17235_/Y _17260_/X VGND VGND VPWR VPWR _17262_/A sky130_fd_sc_hd__or4_4
XANTENNA__15788__A _15795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14472_/Y _14466_/X _14400_/X _14453_/Y VGND VGND VPWR VPWR _25109_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _11685_/A VGND VGND VPWR VPWR _11685_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23078__B2 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16212_ _16217_/A VGND VGND VPWR VPWR _16212_/X sky130_fd_sc_hd__buf_2
X_19000_ _19000_/A VGND VGND VPWR VPWR _19000_/Y sky130_fd_sc_hd__inv_2
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13424_ _13392_/A _23622_/Q VGND VGND VPWR VPWR _13424_/X sky130_fd_sc_hd__or2_4
XFILLER_35_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17192_ _17192_/A VGND VGND VPWR VPWR _17254_/C sky130_fd_sc_hd__inv_2
XANTENNA__22825__B2 _22280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16143_ HWDATA[9] VGND VGND VPWR VPWR _16143_/X sky130_fd_sc_hd__buf_2
X_13355_ _13387_/A _19299_/A VGND VGND VPWR VPWR _13355_/X sky130_fd_sc_hd__or2_4
XFILLER_128_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ _25348_/Q VGND VGND VPWR VPWR _12306_/Y sky130_fd_sc_hd__inv_2
X_16074_ _16073_/Y _15996_/X _15840_/X _15996_/X VGND VGND VPWR VPWR _24704_/D sky130_fd_sc_hd__a2bb2o_4
X_13286_ _13246_/X _23634_/Q VGND VGND VPWR VPWR _13286_/X sky130_fd_sc_hd__or2_4
XFILLER_68_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15025_ _15025_/A VGND VGND VPWR VPWR _15025_/Y sky130_fd_sc_hd__inv_2
X_19902_ _19902_/A VGND VGND VPWR VPWR _19902_/X sky130_fd_sc_hd__buf_2
XANTENNA__24053__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12237_ _25434_/Q VGND VGND VPWR VPWR _12238_/A sky130_fd_sc_hd__inv_2
XFILLER_107_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23250__A1 _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_44_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_89_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21261__B1 _21260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19833_ _19833_/A VGND VGND VPWR VPWR _21745_/B sky130_fd_sc_hd__inv_2
X_12168_ _12167_/X VGND VGND VPWR VPWR _12168_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19764_ _19763_/Y _19759_/X _19740_/X _19759_/X VGND VGND VPWR VPWR _19764_/X sky130_fd_sc_hd__a2bb2o_4
X_12099_ _16183_/A _12054_/X VGND VGND VPWR VPWR _12100_/D sky130_fd_sc_hd__or2_4
X_16976_ _24384_/Q VGND VGND VPWR VPWR _16976_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25259__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18715_ _18705_/B _18704_/X _18707_/X _18712_/B VGND VGND VPWR VPWR _18715_/X sky130_fd_sc_hd__a211o_4
X_15927_ _15845_/A VGND VGND VPWR VPWR _15927_/X sky130_fd_sc_hd__buf_2
X_19695_ _19694_/Y _19690_/X _19599_/X _19690_/X VGND VGND VPWR VPWR _19695_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13771__A _24936_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18646_ _16590_/Y _24126_/Q _16590_/Y _24126_/Q VGND VGND VPWR VPWR _18646_/X sky130_fd_sc_hd__a2bb2o_4
X_15858_ _15852_/A VGND VGND VPWR VPWR _21071_/A sky130_fd_sc_hd__buf_2
XFILLER_64_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16440__B1 _16359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14809_ _14809_/A VGND VGND VPWR VPWR _14810_/A sky130_fd_sc_hd__inv_2
X_18577_ _18393_/Y _18562_/B VGND VGND VPWR VPWR _18577_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12387__A _25451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15789_ _22123_/A VGND VGND VPWR VPWR _21025_/A sky130_fd_sc_hd__buf_2
XFILLER_75_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17528_ _24283_/Q VGND VGND VPWR VPWR _17528_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24894__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17459_ _24194_/Q VGND VGND VPWR VPWR _17459_/X sky130_fd_sc_hd__buf_2
XANTENNA__18074__A _17990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24823__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20470_ _14278_/A _20485_/B _20515_/B VGND VGND VPWR VPWR _20517_/A sky130_fd_sc_hd__and3_4
X_19129_ _19129_/A VGND VGND VPWR VPWR _19130_/A sky130_fd_sc_hd__inv_2
XANTENNA__19693__B1 _19547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14107__A _14381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22140_ _24708_/Q _22135_/X _21024_/A _22139_/X VGND VGND VPWR VPWR _22140_/X sky130_fd_sc_hd__a211o_4
XFILLER_69_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22071_ _22070_/X _22071_/B VGND VGND VPWR VPWR _22071_/X sky130_fd_sc_hd__or2_4
XFILLER_133_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17418__A _16057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16322__A _24615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21022_ _21015_/A VGND VGND VPWR VPWR _21826_/A sky130_fd_sc_hd__inv_2
XFILLER_0_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16274__A3 _16270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_1_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__19748__B2 _19729_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22973_ _22770_/X _22971_/X _22479_/X _24724_/Q _22972_/X VGND VGND VPWR VPWR _22973_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_110_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24712_ _24712_/CLK _16053_/X HRESETn VGND VGND VPWR VPWR _24712_/Q sky130_fd_sc_hd__dfrtp_4
X_21924_ _18307_/X VGND VGND VPWR VPWR _22009_/A sky130_fd_sc_hd__buf_2
XFILLER_55_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16431__B1 _16147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24643_ _24643_/CLK _16248_/X HRESETn VGND VGND VPWR VPWR _24643_/Q sky130_fd_sc_hd__dfrtp_4
X_21855_ _16723_/A VGND VGND VPWR VPWR _23085_/A sky130_fd_sc_hd__buf_2
XANTENNA__16982__A1 _24732_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18708__C1 _18707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _20680_/X _20805_/X _15565_/A _20725_/X VGND VGND VPWR VPWR _20806_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24574_ _24572_/CLK _16432_/X HRESETn VGND VGND VPWR VPWR _15105_/A sky130_fd_sc_hd__dfrtp_4
X_21786_ _21484_/A _21786_/B VGND VGND VPWR VPWR _21786_/X sky130_fd_sc_hd__or2_4
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23525_ _24309_/CLK _20020_/X VGND VGND VPWR VPWR _23525_/Q sky130_fd_sc_hd__dfxtp_4
X_20737_ _20721_/X _20736_/X _15604_/A _20726_/X VGND VGND VPWR VPWR _20737_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18840__A1_N _24561_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24564__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23456_ _23453_/CLK _20201_/X VGND VGND VPWR VPWR _20200_/A sky130_fd_sc_hd__dfxtp_4
X_20668_ _20664_/A _14282_/X VGND VGND VPWR VPWR _20668_/X sky130_fd_sc_hd__or2_4
XFILLER_51_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22407_ _22407_/A _22407_/B VGND VGND VPWR VPWR _22407_/X sky130_fd_sc_hd__and2_4
XFILLER_125_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23387_ _24219_/CLK _23387_/D VGND VGND VPWR VPWR _22390_/A sky130_fd_sc_hd__dfxtp_4
X_20599_ _20447_/X _20455_/B _14089_/X VGND VGND VPWR VPWR _23952_/D sky130_fd_sc_hd__o21a_4
XFILLER_100_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18712__A _24142_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13140_ _13140_/A _13139_/Y VGND VGND VPWR VPWR _13140_/X sky130_fd_sc_hd__and2_4
X_25126_ _24364_/CLK _25126_/D HRESETn VGND VGND VPWR VPWR _25126_/Q sky130_fd_sc_hd__dfstp_4
X_22338_ _22334_/X _22337_/X _18298_/X VGND VGND VPWR VPWR _22338_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_100_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18855__A1_N _24540_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13856__A _23989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13071_ _13002_/B _13071_/B VGND VGND VPWR VPWR _13071_/X sky130_fd_sc_hd__or2_4
XANTENNA__19436__B1 _19389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25057_ _25054_/CLK _14709_/Y HRESETn VGND VGND VPWR VPWR _25057_/Q sky130_fd_sc_hd__dfstp_4
X_22269_ _22265_/X _22267_/X _21290_/C _12296_/A _22268_/X VGND VGND VPWR VPWR _22269_/X
+ sky130_fd_sc_hd__a32o_4
X_12022_ _12020_/A _12021_/A _12020_/Y _12021_/Y VGND VGND VPWR VPWR _12026_/C sky130_fd_sc_hd__o22a_4
X_24008_ _24041_/CLK _24008_/D HRESETn VGND VGND VPWR VPWR _20728_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22888__B _22884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16830_ _16840_/A VGND VGND VPWR VPWR _16830_/X sky130_fd_sc_hd__buf_2
XFILLER_120_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25352__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13973_ _20490_/A _13973_/B VGND VGND VPWR VPWR _25230_/D sky130_fd_sc_hd__or2_4
X_16761_ _24448_/Q VGND VGND VPWR VPWR _16761_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18500_ _18500_/A VGND VGND VPWR VPWR _24173_/D sky130_fd_sc_hd__inv_2
X_12924_ _12924_/A _12902_/X VGND VGND VPWR VPWR _12927_/B sky130_fd_sc_hd__or2_4
X_15712_ _15548_/X _15705_/X _15553_/X _24873_/Q _15711_/X VGND VGND VPWR VPWR _15712_/X
+ sky130_fd_sc_hd__a32o_4
X_16692_ _24477_/Q VGND VGND VPWR VPWR _22598_/A sky130_fd_sc_hd__inv_2
X_19480_ _19480_/A VGND VGND VPWR VPWR _21807_/B sky130_fd_sc_hd__inv_2
XFILLER_111_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16422__B1 _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18431_ _18431_/A _18428_/X _18429_/X _18431_/D VGND VGND VPWR VPWR _18450_/A sky130_fd_sc_hd__or4_4
XFILLER_111_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12855_ _12880_/A _12877_/B VGND VGND VPWR VPWR _12855_/X sky130_fd_sc_hd__or2_4
X_15643_ _16640_/B VGND VGND VPWR VPWR _15643_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17998__A _17990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16973__A1 _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11806_ _11802_/Y _11795_/X _11804_/X _11805_/X VGND VGND VPWR VPWR _11806_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15574_ _24905_/Q VGND VGND VPWR VPWR _15574_/Y sky130_fd_sc_hd__inv_2
X_18362_ _18358_/Y _18361_/Y _18358_/A _18361_/A VGND VGND VPWR VPWR _24189_/D sky130_fd_sc_hd__o22a_4
X_12786_ _12954_/A _24781_/Q _12955_/A _12785_/Y VGND VGND VPWR VPWR _12790_/C sky130_fd_sc_hd__o22a_4
XPHY_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22409__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14521_/X _14524_/X _14483_/A _14517_/X VGND VGND VPWR VPWR _14525_/X sky130_fd_sc_hd__o22a_4
X_17313_ _17252_/C _17311_/A VGND VGND VPWR VPWR _17313_/X sky130_fd_sc_hd__or2_4
XANTENNA__21313__A _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11737_ _21582_/B VGND VGND VPWR VPWR _21066_/A sky130_fd_sc_hd__buf_2
XPHY_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _21194_/A _18293_/B VGND VGND VPWR VPWR _18301_/B sky130_fd_sc_hd__and2_4
XANTENNA__12935__A _22660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22128__B _15708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _20529_/A VGND VGND VPWR VPWR _14456_/Y sky130_fd_sc_hd__inv_2
X_17244_ _24331_/Q VGND VGND VPWR VPWR _17244_/Y sky130_fd_sc_hd__inv_2
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ _13718_/A _24220_/Q _13718_/A _24220_/Q VGND VGND VPWR VPWR _11668_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _13173_/X _13403_/X _13406_/X VGND VGND VPWR VPWR _13407_/X sky130_fd_sc_hd__or3_4
X_17175_ _17246_/C VGND VGND VPWR VPWR _17350_/C sky130_fd_sc_hd__buf_2
XANTENNA__12211__A1 _25427_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24234__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14387_ _14386_/Y _14382_/X _13837_/X _14384_/X VGND VGND VPWR VPWR _25139_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16126_ _16125_/X VGND VGND VPWR VPWR _16126_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16489__B1 _16403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13338_ _13402_/A _13338_/B VGND VGND VPWR VPWR _13338_/X sky130_fd_sc_hd__or2_4
XANTENNA__17686__C1 _17601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16057_ _16057_/A VGND VGND VPWR VPWR _16057_/X sky130_fd_sc_hd__buf_2
X_13269_ _13269_/A _23376_/Q VGND VGND VPWR VPWR _13271_/B sky130_fd_sc_hd__or2_4
XANTENNA__19427__B1 _19426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15008_ _24441_/Q VGND VGND VPWR VPWR _15008_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22982__B1 _25376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19816_ _19814_/Y _19815_/X _19721_/X _19815_/X VGND VGND VPWR VPWR _19816_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22978__A2_N _22974_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25093__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_131_0_HCLK clkbuf_7_65_0_HCLK/X VGND VGND VPWR VPWR _23798_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16661__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19747_ _19747_/A VGND VGND VPWR VPWR _19747_/Y sky130_fd_sc_hd__inv_2
X_16959_ _15990_/Y _24391_/Q _15990_/Y _24391_/Q VGND VGND VPWR VPWR _16959_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_194_0_HCLK clkbuf_7_97_0_HCLK/X VGND VGND VPWR VPWR _24700_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18069__A _18217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22734__B1 _22527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21537__B2 _23100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25022__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19678_ _19678_/A VGND VGND VPWR VPWR _19678_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21207__B _21197_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18402__B2 _18503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18629_ _24531_/Q _24142_/Q _16549_/Y _18705_/A VGND VGND VPWR VPWR _18635_/B sky130_fd_sc_hd__o22a_4
XFILLER_129_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21640_ _21636_/X _21639_/X _13802_/A _18261_/A VGND VGND VPWR VPWR _21640_/X sky130_fd_sc_hd__o22a_4
XFILLER_127_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11789__B1 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21571_ _15010_/Y _22835_/A VGND VGND VPWR VPWR _21571_/X sky130_fd_sc_hd__and2_4
XANTENNA__12450__A1 _12440_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23310_ _23310_/A _23310_/B VGND VGND VPWR VPWR _23310_/X sky130_fd_sc_hd__or2_4
X_20522_ _14279_/A _24066_/Q _20474_/B VGND VGND VPWR VPWR _20522_/X sky130_fd_sc_hd__and3_4
XFILLER_119_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24290_ _24290_/CLK _17660_/Y HRESETn VGND VGND VPWR VPWR _17571_/A sky130_fd_sc_hd__dfrtp_4
X_23241_ _23222_/X _23225_/X _23229_/Y _23240_/X VGND VGND VPWR VPWR HRDATA[28] sky130_fd_sc_hd__a211o_4
X_20453_ _20453_/A _20452_/X VGND VGND VPWR VPWR _20458_/B sky130_fd_sc_hd__and2_4
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23172_ _22798_/A VGND VGND VPWR VPWR _23172_/X sky130_fd_sc_hd__buf_2
X_20384_ _20383_/X _20379_/X _11838_/A _23386_/Q _20381_/X VGND VGND VPWR VPWR _20384_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_106_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22054__A _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22123_ _22123_/A VGND VGND VPWR VPWR _22836_/B sky130_fd_sc_hd__buf_2
XANTENNA__19418__B1 _19349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16052__A _16060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23957__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22054_ _22050_/X _19782_/Y VGND VGND VPWR VPWR _22054_/X sky130_fd_sc_hd__or2_4
XFILLER_43_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22973__B1 _24724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21005_ _21005_/A _21005_/B VGND VGND VPWR VPWR _21005_/X sky130_fd_sc_hd__and2_4
Xclkbuf_7_90_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_90_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16652__B1 _16384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21117__B _11726_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22956_ _12822_/Y _22707_/X _22843_/X _12584_/Y _22844_/X VGND VGND VPWR VPWR _22956_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__16404__B1 _16403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21907_ _21904_/A _20088_/Y VGND VGND VPWR VPWR _21907_/X sky130_fd_sc_hd__or2_4
XFILLER_28_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22887_ _14913_/A _22523_/A _22524_/A _22886_/X VGND VGND VPWR VPWR _22888_/C sky130_fd_sc_hd__a211o_4
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20751__A2 _20745_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12640_ _12622_/A _12638_/X _12648_/A _12635_/B VGND VGND VPWR VPWR _12641_/A sky130_fd_sc_hd__a211o_4
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24626_ _24330_/CLK _16294_/X HRESETn VGND VGND VPWR VPWR _24626_/Q sky130_fd_sc_hd__dfrtp_4
X_21838_ _24506_/Q _21312_/X _22997_/A _21837_/X VGND VGND VPWR VPWR _21839_/C sky130_fd_sc_hd__a211o_4
XFILLER_43_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24745__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ _12570_/Y _24855_/Q _12570_/Y _24855_/Q VGND VGND VPWR VPWR _12578_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12441__A1 _12286_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24557_ _24557_/CLK _16482_/X HRESETn VGND VGND VPWR VPWR _24557_/Q sky130_fd_sc_hd__dfrtp_4
X_21769_ _21596_/A _21769_/B VGND VGND VPWR VPWR _21769_/X sky130_fd_sc_hd__or2_4
XANTENNA__12755__A _22546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ _25164_/Q _14302_/X _25163_/Q _14307_/X VGND VGND VPWR VPWR _14310_/X sky130_fd_sc_hd__o22a_4
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23508_ _24187_/CLK _20067_/X VGND VGND VPWR VPWR _23508_/Q sky130_fd_sc_hd__dfxtp_4
X_15290_ _24465_/Q VGND VGND VPWR VPWR _15387_/B sky130_fd_sc_hd__inv_2
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24488_ _24487_/CLK _24488_/D HRESETn VGND VGND VPWR VPWR _24488_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14241_ _25181_/Q VGND VGND VPWR VPWR _14241_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23439_ _23904_/CLK _23439_/D VGND VGND VPWR VPWR _13373_/B sky130_fd_sc_hd__dfxtp_4
X_14172_ _14171_/X VGND VGND VPWR VPWR _14173_/B sky130_fd_sc_hd__buf_2
X_13123_ _13121_/Y _13123_/B VGND VGND VPWR VPWR _13123_/X sky130_fd_sc_hd__and2_4
XFILLER_124_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25109_ _23959_/CLK _25109_/D HRESETn VGND VGND VPWR VPWR _25109_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19409__B1 _19407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15143__B1 _24973_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18980_ _18980_/A VGND VGND VPWR VPWR _18980_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25533__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13054_ _13054_/A _13061_/A _13057_/A _13067_/B VGND VGND VPWR VPWR _13060_/B sky130_fd_sc_hd__or4_4
X_17931_ _17957_/A _17931_/B _17931_/C VGND VGND VPWR VPWR _17931_/X sky130_fd_sc_hd__and3_4
X_12005_ _24087_/Q _11992_/B _12004_/Y VGND VGND VPWR VPWR _12006_/A sky130_fd_sc_hd__o21a_4
X_17862_ _16918_/Y _17862_/B VGND VGND VPWR VPWR _17863_/C sky130_fd_sc_hd__or2_4
XFILLER_120_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18632__B2 _18792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19601_ _23671_/Q VGND VGND VPWR VPWR _19601_/Y sky130_fd_sc_hd__inv_2
X_16813_ _24424_/Q VGND VGND VPWR VPWR _16813_/Y sky130_fd_sc_hd__inv_2
X_17793_ _17741_/Y _17792_/X VGND VGND VPWR VPWR _17794_/B sky130_fd_sc_hd__or2_4
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_204_0_HCLK clkbuf_8_205_0_HCLK/A VGND VGND VPWR VPWR _24840_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22130__C _22130_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19532_ _19532_/A VGND VGND VPWR VPWR _21174_/B sky130_fd_sc_hd__inv_2
X_16744_ _15042_/Y _16739_/X _16393_/X _16743_/X VGND VGND VPWR VPWR _24457_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21027__B _21027_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13956_ _13956_/A VGND VGND VPWR VPWR _13958_/A sky130_fd_sc_hd__inv_2
XANTENNA__14210__A _20657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12907_ _25376_/Q _12906_/Y VGND VGND VPWR VPWR _12907_/X sky130_fd_sc_hd__or2_4
X_19463_ _19461_/Y _19459_/X _19462_/X _19459_/X VGND VGND VPWR VPWR _19463_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13887_ _13927_/B VGND VGND VPWR VPWR _13893_/B sky130_fd_sc_hd__buf_2
X_16675_ _24484_/Q VGND VGND VPWR VPWR _22872_/A sky130_fd_sc_hd__inv_2
XANTENNA__16946__B2 _16927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18414_ _18414_/A VGND VGND VPWR VPWR _18481_/B sky130_fd_sc_hd__inv_2
X_12838_ _12838_/A VGND VGND VPWR VPWR _12979_/A sky130_fd_sc_hd__buf_2
X_15626_ _15561_/X VGND VGND VPWR VPWR _15626_/X sky130_fd_sc_hd__buf_2
XANTENNA__24486__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19394_ _18165_/B VGND VGND VPWR VPWR _19394_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22139__A _15708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21043__A _11720_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18345_ _18345_/A VGND VGND VPWR VPWR _18345_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24415__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12769_ _24780_/Q VGND VGND VPWR VPWR _12769_/Y sky130_fd_sc_hd__inv_2
X_15557_ _16640_/A _15777_/A VGND VGND VPWR VPWR _15560_/A sky130_fd_sc_hd__or2_4
XANTENNA__12665__A _12665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14508_ _14503_/B VGND VGND VPWR VPWR _14508_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_2_1_0_HCLK_A clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15488_ _15487_/X VGND VGND VPWR VPWR _24064_/D sky130_fd_sc_hd__buf_2
X_18276_ _17708_/A VGND VGND VPWR VPWR _20000_/C sky130_fd_sc_hd__buf_2
XANTENNA__12384__B _13008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20891__A1_N _20882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17227_ _24627_/Q _17234_/A _16354_/Y _24332_/Q VGND VGND VPWR VPWR _17229_/C sky130_fd_sc_hd__a2bb2o_4
X_14439_ _25123_/Q VGND VGND VPWR VPWR _14439_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21697__B _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17659__C1 _17590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17158_ _17156_/Y _17157_/X _17160_/C VGND VGND VPWR VPWR _24363_/D sky130_fd_sc_hd__and3_4
X_16109_ _16108_/Y _16106_/X _11771_/X _16106_/X VGND VGND VPWR VPWR _24691_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17089_ _17089_/A VGND VGND VPWR VPWR _17089_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25274__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_14_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__25203__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19820__B1 _19771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16600__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22810_ _22836_/B VGND VGND VPWR VPWR _22810_/X sky130_fd_sc_hd__buf_2
XFILLER_38_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23790_ _23846_/CLK _23790_/D VGND VGND VPWR VPWR _19258_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_84_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18387__B1 _24178_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12120__B1 _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13463__A3 _13462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22741_ _22476_/X _22740_/X _21285_/A _24822_/Q _22480_/X VGND VGND VPWR VPWR _22741_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_1_0_1_HCLK clkbuf_1_0_1_HCLK/A VGND VGND VPWR VPWR clkbuf_2_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25460_ _25461_/CLK _12115_/X HRESETn VGND VGND VPWR VPWR _12113_/A sky130_fd_sc_hd__dfrtp_4
X_22672_ _20734_/Y _22988_/A _20873_/Y _21588_/X VGND VGND VPWR VPWR _22672_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24411_ _24407_/CLK _24411_/D HRESETn VGND VGND VPWR VPWR _14900_/A sky130_fd_sc_hd__dfrtp_4
X_21623_ _21623_/A _20181_/Y VGND VGND VPWR VPWR _21624_/C sky130_fd_sc_hd__or2_4
XANTENNA__24156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25391_ _25411_/CLK _25391_/D HRESETn VGND VGND VPWR VPWR _12590_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16047__A _16060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24342_ _24345_/CLK _24342_/D HRESETn VGND VGND VPWR VPWR _22702_/A sky130_fd_sc_hd__dfrtp_4
X_21554_ _21554_/A VGND VGND VPWR VPWR _21554_/Y sky130_fd_sc_hd__inv_2
X_20505_ _14278_/A _20474_/B _20505_/C VGND VGND VPWR VPWR _20517_/D sky130_fd_sc_hd__and3_4
XANTENNA__15886__A _15713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23156__A1_N _12290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24273_ _24682_/CLK _17782_/Y HRESETn VGND VGND VPWR VPWR _24273_/Q sky130_fd_sc_hd__dfrtp_4
X_21485_ _21485_/A _21485_/B _21484_/X VGND VGND VPWR VPWR _21485_/X sky130_fd_sc_hd__and3_4
XFILLER_14_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23224_ _17261_/B _22475_/X _25383_/Q _22435_/X VGND VGND VPWR VPWR _23224_/X sky130_fd_sc_hd__a2bb2o_4
X_20436_ _20428_/B _20427_/C _20433_/X VGND VGND VPWR VPWR _20436_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23155_ _23114_/A _23155_/B _23155_/C _23154_/X VGND VGND VPWR VPWR _23155_/X sky130_fd_sc_hd__or4_4
X_20367_ _22027_/B _20361_/X _19618_/A _20366_/X VGND VGND VPWR VPWR _23393_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22106_ _12278_/B _15784_/B _16928_/Y _22821_/A VGND VGND VPWR VPWR _22106_/X sky130_fd_sc_hd__o22a_4
XFILLER_121_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23086_ _22819_/X _23077_/Y _23081_/Y _23085_/X VGND VGND VPWR VPWR _23094_/C sky130_fd_sc_hd__a211o_4
X_20298_ _20298_/A VGND VGND VPWR VPWR _20298_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22037_ _22036_/A _19604_/Y VGND VGND VPWR VPWR _22037_/X sky130_fd_sc_hd__or2_4
XFILLER_0_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19811__B1 _19715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24997__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13810_ _16720_/A VGND VGND VPWR VPWR _13810_/X sky130_fd_sc_hd__buf_2
XFILLER_29_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14790_ _18079_/A _14789_/Y _13630_/A _14659_/B VGND VGND VPWR VPWR _14790_/X sky130_fd_sc_hd__o22a_4
XFILLER_75_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24926__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23988_ _25043_/CLK _23988_/D HRESETn VGND VGND VPWR VPWR _14870_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_21_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13741_ _13741_/A _16630_/A _13741_/C VGND VGND VPWR VPWR _13742_/A sky130_fd_sc_hd__and3_4
XFILLER_84_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22939_ _22939_/A _21048_/B VGND VGND VPWR VPWR _22939_/X sky130_fd_sc_hd__or2_4
XFILLER_21_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_34_0_HCLK clkbuf_8_34_0_HCLK/A VGND VGND VPWR VPWR _23826_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_5_18_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13672_ _25286_/Q _13670_/X _13671_/Y VGND VGND VPWR VPWR _25286_/D sky130_fd_sc_hd__o21a_4
X_16460_ _16466_/A VGND VGND VPWR VPWR _16461_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_97_0_HCLK clkbuf_7_48_0_HCLK/X VGND VGND VPWR VPWR _23959_/CLK sky130_fd_sc_hd__clkbuf_1
X_12623_ _12623_/A _12693_/A _12623_/C VGND VGND VPWR VPWR _12626_/B sky130_fd_sc_hd__or3_4
X_15411_ _15390_/X _15411_/B _15407_/X VGND VGND VPWR VPWR _15411_/X sky130_fd_sc_hd__and3_4
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16391_ _24592_/Q VGND VGND VPWR VPWR _16391_/Y sky130_fd_sc_hd__inv_2
X_24609_ _24889_/CLK _16341_/X HRESETn VGND VGND VPWR VPWR _24609_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15342_ _15338_/A _15338_/B VGND VGND VPWR VPWR _15343_/C sky130_fd_sc_hd__nand2_4
X_18130_ _15695_/X _18114_/X _18129_/X _24233_/Q _18019_/X VGND VGND VPWR VPWR _18130_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ _25406_/Q VGND VGND VPWR VPWR _12681_/A sky130_fd_sc_hd__inv_2
XFILLER_106_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15273_ _25000_/Q _15272_/Y VGND VGND VPWR VPWR _15273_/X sky130_fd_sc_hd__or2_4
X_18061_ _17963_/X _18060_/X _24234_/Q _18021_/X VGND VGND VPWR VPWR _24234_/D sky130_fd_sc_hd__o22a_4
X_12485_ _12203_/X _12471_/X _12412_/A _12481_/Y VGND VGND VPWR VPWR _12485_/X sky130_fd_sc_hd__a211o_4
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12178__B1 _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14224_ _14224_/A VGND VGND VPWR VPWR _14224_/X sky130_fd_sc_hd__buf_2
X_17012_ _16069_/Y _17039_/A _24704_/Q _16993_/Y VGND VGND VPWR VPWR _17016_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22406__B _22406_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14155_ _14146_/X _14154_/Y _25124_/Q _14146_/X VGND VGND VPWR VPWR _25204_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11829__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12817__A1_N _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13106_ _13106_/A _13113_/A VGND VGND VPWR VPWR _13106_/X sky130_fd_sc_hd__or2_4
X_14086_ _23995_/Q _14078_/A _14073_/X _13982_/A _14084_/X VGND VGND VPWR VPWR _14086_/X
+ sky130_fd_sc_hd__a32o_4
X_18963_ _13409_/B VGND VGND VPWR VPWR _18963_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22422__A _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13037_ _25345_/Q _13037_/B VGND VGND VPWR VPWR _13037_/X sky130_fd_sc_hd__or2_4
X_17914_ _15915_/B _17920_/C VGND VGND VPWR VPWR _17914_/Y sky130_fd_sc_hd__nor2_4
X_18894_ _20984_/A VGND VGND VPWR VPWR _18894_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17845_ _17737_/X VGND VGND VPWR VPWR _17874_/A sky130_fd_sc_hd__buf_2
XFILLER_66_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24667__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17776_ _17776_/A VGND VGND VPWR VPWR _17776_/Y sky130_fd_sc_hd__inv_2
X_14988_ _15219_/A _24451_/Q _15219_/A _24451_/Q VGND VGND VPWR VPWR _14996_/A sky130_fd_sc_hd__a2bb2o_4
X_19515_ _19515_/A VGND VGND VPWR VPWR _19528_/A sky130_fd_sc_hd__inv_2
X_16727_ _24464_/Q VGND VGND VPWR VPWR _16727_/Y sky130_fd_sc_hd__inv_2
X_13939_ _13956_/A _13939_/B _13930_/D _13958_/D VGND VGND VPWR VPWR _13939_/X sky130_fd_sc_hd__or4_4
XANTENNA__20176__B1 _20085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19446_ _19445_/X VGND VGND VPWR VPWR _19446_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16658_ _16658_/A VGND VGND VPWR VPWR _16658_/X sky130_fd_sc_hd__buf_2
XFILLER_34_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15609_ _24891_/Q VGND VGND VPWR VPWR _15609_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_5_5_0_HCLK clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19377_ _19014_/A _19038_/B _19038_/C _19038_/D VGND VGND VPWR VPWR _19377_/X sky130_fd_sc_hd__and4_4
X_16589_ _16587_/Y _16583_/X _16231_/X _16588_/X VGND VGND VPWR VPWR _24516_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18328_ _17466_/Y _19219_/C _17467_/Y VGND VGND VPWR VPWR _19683_/C sky130_fd_sc_hd__or3_4
XFILLER_50_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21501__A _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18259_ _18259_/A VGND VGND VPWR VPWR _18259_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25455__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21270_ _22505_/A VGND VGND VPWR VPWR _21270_/X sky130_fd_sc_hd__buf_2
XFILLER_116_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12842__B _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20221_ _20221_/A VGND VGND VPWR VPWR _20221_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20152_ _22197_/B _20149_/X _20082_/X _20149_/X VGND VGND VPWR VPWR _23475_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22332__A _21944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24960_ _24957_/CLK _15440_/X HRESETn VGND VGND VPWR VPWR _13924_/A sky130_fd_sc_hd__dfrtp_4
X_20083_ _22194_/B _20078_/X _20082_/X _20078_/X VGND VGND VPWR VPWR _23499_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16607__B1 _16521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23911_ _23846_/CLK _23911_/D VGND VGND VPWR VPWR _23911_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24891_ _24893_/CLK _24891_/D HRESETn VGND VGND VPWR VPWR _24891_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17280__B1 _17279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23842_ _23854_/CLK _19113_/X VGND VGND VPWR VPWR _13263_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22156__A1 _16608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12289__B _12252_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24337__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_250_0_HCLK clkbuf_7_125_0_HCLK/X VGND VGND VPWR VPWR _23370_/CLK sky130_fd_sc_hd__clkbuf_1
X_23773_ _23618_/CLK _19308_/X VGND VGND VPWR VPWR _13451_/B sky130_fd_sc_hd__dfxtp_4
X_20985_ _20479_/A _23956_/Q _20490_/A VGND VGND VPWR VPWR _23956_/D sky130_fd_sc_hd__a21o_4
XANTENNA__13841__B1 _13840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25512_ _25514_/CLK _11843_/X HRESETn VGND VGND VPWR VPWR _25512_/Q sky130_fd_sc_hd__dfrtp_4
X_22724_ _24416_/Q _22523_/X _22524_/X _22723_/X VGND VGND VPWR VPWR _22725_/C sky130_fd_sc_hd__a211o_4
XFILLER_41_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25443_ _25449_/CLK _12425_/X HRESETn VGND VGND VPWR VPWR _25443_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15594__B1 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22655_ _22655_/A _22654_/X VGND VGND VPWR VPWR _22655_/X sky130_fd_sc_hd__or2_4
XFILLER_55_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21606_ _21599_/X _21605_/X _14712_/X VGND VGND VPWR VPWR _21606_/X sky130_fd_sc_hd__o21a_4
X_25374_ _25374_/CLK _25374_/D HRESETn VGND VGND VPWR VPWR _12778_/A sky130_fd_sc_hd__dfrtp_4
X_22586_ _22736_/A _22583_/X _22586_/C VGND VGND VPWR VPWR _22586_/X sky130_fd_sc_hd__and3_4
XANTENNA__21411__A _23100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24325_ _23964_/CLK _24325_/D HRESETn VGND VGND VPWR VPWR _20992_/B sky130_fd_sc_hd__dfstp_4
X_21537_ _17199_/Y _21303_/X _25357_/Q _23100_/A VGND VGND VPWR VPWR _21538_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23972__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25196__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12270_ _12269_/Y _22267_/A _12264_/X _24738_/Q VGND VGND VPWR VPWR _12271_/D sky130_fd_sc_hd__a2bb2o_4
X_24256_ _24673_/CLK _24256_/D HRESETn VGND VGND VPWR VPWR _17744_/A sky130_fd_sc_hd__dfrtp_4
X_21468_ _21464_/X _21467_/X _18299_/X VGND VGND VPWR VPWR _21468_/X sky130_fd_sc_hd__o21a_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15543__A2_N _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23207_ _23207_/A _23204_/X _23207_/C VGND VGND VPWR VPWR _23208_/D sky130_fd_sc_hd__and3_4
X_20419_ _24063_/D _20419_/B VGND VGND VPWR VPWR _20419_/X sky130_fd_sc_hd__or2_4
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22092__B1 _22090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18835__A1 _24563_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24187_ _24187_/CLK _18366_/X HRESETn VGND VGND VPWR VPWR _24187_/Q sky130_fd_sc_hd__dfrtp_4
X_21399_ _21381_/A _20142_/Y VGND VGND VPWR VPWR _21399_/X sky130_fd_sc_hd__or2_4
XANTENNA__18835__B2 _18705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12471__C _12278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23983__D scl_i_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16846__B1 _16528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23138_ _23208_/A _23128_/Y _23133_/X _23138_/D VGND VGND VPWR VPWR _23138_/X sky130_fd_sc_hd__or4_4
XFILLER_49_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19535__B _14192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17336__A _17260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15960_ _15938_/X VGND VGND VPWR VPWR _15960_/X sky130_fd_sc_hd__buf_2
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23069_ _24558_/Q _23069_/B _23005_/C VGND VGND VPWR VPWR _23069_/X sky130_fd_sc_hd__and3_4
XFILLER_103_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14911_ _25013_/Q VGND VGND VPWR VPWR _15067_/A sky130_fd_sc_hd__inv_2
XFILLER_118_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15891_ _15886_/X _15887_/X _11803_/X _22708_/A _15888_/X VGND VGND VPWR VPWR _24786_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_60_0_HCLK clkbuf_6_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17630_ _17630_/A _17630_/B VGND VGND VPWR VPWR _17631_/C sky130_fd_sc_hd__or2_4
X_14842_ _14810_/X _14841_/X _25183_/Q _14835_/X VGND VGND VPWR VPWR _14842_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__24760__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17561_ _24301_/Q VGND VGND VPWR VPWR _17612_/A sky130_fd_sc_hd__inv_2
XFILLER_84_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23048__A1_N _12244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24078__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11985_ _11654_/A _11654_/B _11984_/Y VGND VGND VPWR VPWR _11985_/Y sky130_fd_sc_hd__a21oi_4
X_14773_ _14772_/X VGND VGND VPWR VPWR _14776_/B sky130_fd_sc_hd__inv_2
XFILLER_91_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13832__B1 _11825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19300_ _19299_/Y _19295_/X _19232_/X _19295_/X VGND VGND VPWR VPWR _19300_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16512_ _16510_/Y _16511_/X _16242_/X _16511_/X VGND VGND VPWR VPWR _16512_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13724_ _13685_/X _13723_/Y _13721_/X _13714_/X _25273_/Q VGND VGND VPWR VPWR _13724_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24007__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17492_ _11815_/Y _24289_/Q _11815_/Y _24289_/Q VGND VGND VPWR VPWR _17497_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19231_ _13340_/B VGND VGND VPWR VPWR _19231_/Y sky130_fd_sc_hd__inv_2
X_16443_ _15115_/Y _16437_/X _16442_/X _16437_/X VGND VGND VPWR VPWR _24569_/D sky130_fd_sc_hd__a2bb2o_4
X_13655_ _13655_/A _13655_/B VGND VGND VPWR VPWR _13656_/B sky130_fd_sc_hd__or2_4
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _12606_/A VGND VGND VPWR VPWR _12622_/A sky130_fd_sc_hd__inv_2
X_19162_ _19162_/A VGND VGND VPWR VPWR _19162_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13586_ _25242_/Q _14560_/B _13831_/A _14592_/A VGND VGND VPWR VPWR _13587_/D sky130_fd_sc_hd__a2bb2o_4
X_16374_ _16381_/A VGND VGND VPWR VPWR _16375_/A sky130_fd_sc_hd__buf_2
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22417__A _22383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18113_ _18224_/A _18109_/X _18113_/C VGND VGND VPWR VPWR _18113_/X sky130_fd_sc_hd__or3_4
XFILLER_8_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12537_ _25396_/Q _24850_/Q _12707_/A _12536_/Y VGND VGND VPWR VPWR _12537_/X sky130_fd_sc_hd__o22a_4
X_15325_ _15087_/Y _15325_/B _15331_/A _15316_/X VGND VGND VPWR VPWR _15325_/X sky130_fd_sc_hd__or4_4
X_19093_ _23849_/Q VGND VGND VPWR VPWR _21888_/B sky130_fd_sc_hd__inv_2
XFILLER_117_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18044_ _18000_/A _18042_/X _18044_/C VGND VGND VPWR VPWR _18048_/B sky130_fd_sc_hd__and3_4
X_12468_ _12196_/Y _12382_/X VGND VGND VPWR VPWR _12509_/B sky130_fd_sc_hd__or2_4
X_15256_ _15262_/A _15251_/B _15250_/X VGND VGND VPWR VPWR _15256_/X sky130_fd_sc_hd__or3_4
X_14207_ _14207_/A VGND VGND VPWR VPWR _14207_/Y sky130_fd_sc_hd__inv_2
X_15187_ _15187_/A _15185_/A VGND VGND VPWR VPWR _15188_/C sky130_fd_sc_hd__or2_4
X_12399_ _12399_/A _12398_/Y VGND VGND VPWR VPWR _12401_/B sky130_fd_sc_hd__or2_4
XANTENNA__18630__A _18630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14138_ _14125_/X _14137_/Y _14117_/C _14125_/X VGND VGND VPWR VPWR _14138_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19995_ _19995_/A VGND VGND VPWR VPWR _19995_/X sky130_fd_sc_hd__buf_2
XFILLER_67_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13774__A _13593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14069_ _14078_/A VGND VGND VPWR VPWR _14069_/X sky130_fd_sc_hd__buf_2
X_18946_ _18945_/X VGND VGND VPWR VPWR _18946_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24848__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18877_ _23939_/Q _18876_/X VGND VGND VPWR VPWR _20571_/A sky130_fd_sc_hd__or2_4
XFILLER_80_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20936__A2 _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17828_ _17758_/D _17818_/D _17780_/X _17826_/B VGND VGND VPWR VPWR _17829_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24430__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17759_ _17759_/A _17753_/Y _17759_/C _17758_/X VGND VGND VPWR VPWR _17760_/B sky130_fd_sc_hd__or4_4
XANTENNA__13823__B1 _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18077__A _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20770_ _20770_/A VGND VGND VPWR VPWR _20770_/X sky130_fd_sc_hd__buf_2
XFILLER_39_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19429_ _19428_/Y _19425_/X _19404_/X _19425_/X VGND VGND VPWR VPWR _23731_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15576__B1 _11764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_80_0_HCLK clkbuf_8_81_0_HCLK/A VGND VGND VPWR VPWR _23967_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22440_ _22436_/X _22438_/X _22440_/C VGND VGND VPWR VPWR _22440_/X sky130_fd_sc_hd__or3_4
X_22371_ _21618_/A _22371_/B VGND VGND VPWR VPWR _22371_/X sky130_fd_sc_hd__or2_4
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16325__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24110_ _25199_/CLK _18888_/X HRESETn VGND VGND VPWR VPWR _24110_/Q sky130_fd_sc_hd__dfstp_4
X_21322_ _21322_/A _22298_/B VGND VGND VPWR VPWR _21322_/X sky130_fd_sc_hd__or2_4
Xclkbuf_2_0_0_HCLK clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_2_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_25090_ _25137_/CLK _25090_/D HRESETn VGND VGND VPWR VPWR _21334_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24041_ _24041_/CLK _24041_/D HRESETn VGND VGND VPWR VPWR _24041_/Q sky130_fd_sc_hd__dfrtp_4
X_21253_ _21253_/A _20061_/Y VGND VGND VPWR VPWR _21254_/C sky130_fd_sc_hd__or2_4
XFILLER_116_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20204_ _20202_/Y _20203_/X _16879_/A _20203_/X VGND VGND VPWR VPWR _23455_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16828__B1 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21184_ _21184_/A _21184_/B VGND VGND VPWR VPWR _21186_/B sky130_fd_sc_hd__or2_4
XANTENNA__22062__A _14682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20135_ _23481_/Q VGND VGND VPWR VPWR _21906_/B sky130_fd_sc_hd__inv_2
XANTENNA__15500__B1 HADDR[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24589__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16060__A _16060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22997__A _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20066_ _20065_/Y VGND VGND VPWR VPWR _20066_/X sky130_fd_sc_hd__buf_2
XANTENNA__24518__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24943_ _24943_/CLK _15469_/X HRESETn VGND VGND VPWR VPWR _15467_/A sky130_fd_sc_hd__dfstp_4
XFILLER_86_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_4_0_HCLK_A clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24874_ _23818_/CLK _15699_/X HRESETn VGND VGND VPWR VPWR _15681_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23825_ _25264_/CLK _23825_/D VGND VGND VPWR VPWR _19162_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24100__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11770_ _25530_/Q VGND VGND VPWR VPWR _11770_/Y sky130_fd_sc_hd__inv_2
X_23756_ _23772_/CLK _19357_/X VGND VGND VPWR VPWR _17945_/B sky130_fd_sc_hd__dfxtp_4
X_20968_ _20968_/A _14380_/X VGND VGND VPWR VPWR _23921_/D sky130_fd_sc_hd__and2_4
XFILLER_57_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22707_ _23097_/A VGND VGND VPWR VPWR _22707_/X sky130_fd_sc_hd__buf_2
X_23687_ _23689_/CLK _19554_/X VGND VGND VPWR VPWR _23687_/Q sky130_fd_sc_hd__dfxtp_4
X_20899_ _20882_/X _20898_/X _24484_/Q _20886_/X VGND VGND VPWR VPWR _24047_/D sky130_fd_sc_hd__a2bb2o_4
X_13440_ _13440_/A _23371_/Q VGND VGND VPWR VPWR _13440_/X sky130_fd_sc_hd__or2_4
XANTENNA__25377__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_108_0_HCLK clkbuf_7_54_0_HCLK/X VGND VGND VPWR VPWR _24885_/CLK sky130_fd_sc_hd__clkbuf_1
X_25426_ _25385_/CLK _12492_/X HRESETn VGND VGND VPWR VPWR _25426_/Q sky130_fd_sc_hd__dfrtp_4
X_22638_ _22638_/A VGND VGND VPWR VPWR _22638_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25306__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13371_ _13260_/X _13369_/X _13370_/X VGND VGND VPWR VPWR _13371_/X sky130_fd_sc_hd__and3_4
X_25357_ _25356_/CLK _25357_/D HRESETn VGND VGND VPWR VPWR _25357_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20312__B1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22569_ _22568_/X VGND VGND VPWR VPWR _22570_/D sky130_fd_sc_hd__inv_2
XANTENNA__16235__A _11809_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12322_ _25346_/Q _24831_/Q _13030_/A _12321_/Y VGND VGND VPWR VPWR _12326_/C sky130_fd_sc_hd__o22a_4
X_15110_ _15322_/A _24596_/Q _15309_/C _15109_/Y VGND VGND VPWR VPWR _15120_/A sky130_fd_sc_hd__o22a_4
XFILLER_16_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16090_ _23278_/A VGND VGND VPWR VPWR _16090_/Y sky130_fd_sc_hd__inv_2
X_24308_ _24309_/CLK _24308_/D HRESETn VGND VGND VPWR VPWR _24308_/Q sky130_fd_sc_hd__dfrtp_4
X_25288_ _25478_/CLK _13642_/X HRESETn VGND VGND VPWR VPWR _13527_/B sky130_fd_sc_hd__dfstp_4
XFILLER_103_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15041_ _25001_/Q _15028_/Y _14886_/X _24444_/Q VGND VGND VPWR VPWR _15041_/X sky130_fd_sc_hd__a2bb2o_4
X_12253_ _12252_/Y _24757_/Q _25430_/Q _12190_/Y VGND VGND VPWR VPWR _12253_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24239_ _23516_/CLK _17922_/X HRESETn VGND VGND VPWR VPWR _13541_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12184_ _12184_/A VGND VGND VPWR VPWR _12277_/A sky130_fd_sc_hd__inv_2
XFILLER_64_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18800_ _18792_/B _18792_/C _18724_/A _18796_/Y VGND VGND VPWR VPWR _18800_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17492__B1 _11815_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19780_ _19780_/A VGND VGND VPWR VPWR _19780_/X sky130_fd_sc_hd__buf_2
XFILLER_110_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16992_ _24720_/Q _17034_/B _16063_/Y _16994_/A VGND VGND VPWR VPWR _16998_/A sky130_fd_sc_hd__a2bb2o_4
X_18731_ _18674_/Y _18728_/X VGND VGND VPWR VPWR _18731_/X sky130_fd_sc_hd__or2_4
X_15943_ _12255_/Y _15939_/X _15942_/X _15939_/X VGND VGND VPWR VPWR _15943_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24259__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13744__D _13588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18662_ _16547_/Y _18671_/A _16547_/Y _18671_/A VGND VGND VPWR VPWR _18666_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15874_ _15850_/X _15857_/X _15723_/X _24798_/Q _15864_/X VGND VGND VPWR VPWR _15874_/X
+ sky130_fd_sc_hd__a32o_4
X_17613_ _17616_/A _17616_/B VGND VGND VPWR VPWR _17617_/B sky130_fd_sc_hd__or2_4
X_14825_ _14824_/X VGND VGND VPWR VPWR _14825_/X sky130_fd_sc_hd__buf_2
X_18593_ _24146_/Q _18592_/Y VGND VGND VPWR VPWR _18594_/B sky130_fd_sc_hd__or2_4
XFILLER_40_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13805__B1 _13803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11842__A _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17544_ _25529_/Q _17543_/Y _11780_/Y _24298_/Q VGND VGND VPWR VPWR _17545_/D sky130_fd_sc_hd__a2bb2o_4
X_14756_ _21372_/A VGND VGND VPWR VPWR _21385_/A sky130_fd_sc_hd__buf_2
XFILLER_17_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11968_ _11704_/A _11959_/X _11966_/Y _11961_/A _11967_/X VGND VGND VPWR VPWR _11968_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17547__B2 _24308_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13707_ _13721_/A VGND VGND VPWR VPWR _13707_/X sky130_fd_sc_hd__buf_2
X_17475_ _17474_/A VGND VGND VPWR VPWR _17476_/A sky130_fd_sc_hd__inv_2
XFILLER_32_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11899_ _11899_/A VGND VGND VPWR VPWR _11899_/Y sky130_fd_sc_hd__inv_2
X_14687_ _14679_/A VGND VGND VPWR VPWR _21245_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_67_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_67_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19214_ _18190_/B VGND VGND VPWR VPWR _19214_/Y sky130_fd_sc_hd__inv_2
X_16426_ _16433_/A VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__buf_2
XFILLER_38_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13638_ _13638_/A VGND VGND VPWR VPWR _13638_/X sky130_fd_sc_hd__buf_2
XFILLER_32_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13033__A1 _12299_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14230__B1 _13840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25047__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19145_ _19143_/Y _19144_/X _19077_/X _19144_/X VGND VGND VPWR VPWR _19145_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16357_ _16354_/Y _16350_/X _16355_/X _16356_/X VGND VGND VPWR VPWR _24603_/D sky130_fd_sc_hd__a2bb2o_4
X_13569_ _25255_/Q VGND VGND VPWR VPWR _13569_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23967__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15308_ _15087_/Y _15325_/B VGND VGND VPWR VPWR _15308_/X sky130_fd_sc_hd__or2_4
X_19076_ _19062_/Y VGND VGND VPWR VPWR _19076_/X sky130_fd_sc_hd__buf_2
XANTENNA__16996__A1_N _16044_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16288_ _16280_/X VGND VGND VPWR VPWR _16288_/X sky130_fd_sc_hd__buf_2
XANTENNA__12392__B _12385_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18027_ _18023_/X _18027_/B _18026_/X VGND VGND VPWR VPWR _18027_/X sky130_fd_sc_hd__and3_4
X_15239_ _15239_/A _15239_/B VGND VGND VPWR VPWR _15240_/A sky130_fd_sc_hd__or2_4
XANTENNA__15730__B1 _24865_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19472__B2 _19471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19978_ _11928_/A VGND VGND VPWR VPWR _19978_/X sky130_fd_sc_hd__buf_2
XANTENNA__24682__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18929_ _13272_/B VGND VGND VPWR VPWR _18929_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23020__A2 _22833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24611__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_HCLK HCLK VGND VGND VPWR VPWR clkbuf_0_HCLK/X sky130_fd_sc_hd__clkbuf_16
X_21940_ _21936_/X _21939_/X _17722_/A VGND VGND VPWR VPWR _21940_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19191__A _19055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23308__B1 _24734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18983__B1 _18940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21871_ _22287_/A _21865_/X _22962_/A _21870_/X VGND VGND VPWR VPWR _21875_/A sky130_fd_sc_hd__a211o_4
XANTENNA__12848__A _25376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23610_ _23609_/CLK _23610_/D VGND VGND VPWR VPWR _23610_/Q sky130_fd_sc_hd__dfxtp_4
X_20822_ _16716_/Y _20815_/X _20818_/X _20821_/Y VGND VGND VPWR VPWR _20823_/A sky130_fd_sc_hd__o22a_4
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24590_ _24995_/CLK _16397_/X HRESETn VGND VGND VPWR VPWR _24590_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23541_ _24309_/CLK _19969_/X VGND VGND VPWR VPWR _19968_/A sky130_fd_sc_hd__dfxtp_4
X_20753_ _13119_/A VGND VGND VPWR VPWR _20754_/C sky130_fd_sc_hd__inv_2
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12286__C _12286_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25470__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23472_ _23496_/CLK _23472_/D VGND VGND VPWR VPWR _23472_/Q sky130_fd_sc_hd__dfxtp_4
X_20684_ _15636_/Y _20677_/X _20680_/X _20683_/Y VGND VGND VPWR VPWR _20685_/A sky130_fd_sc_hd__o22a_4
XANTENNA__23087__A2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25211_ _25093_/CLK _25211_/D HRESETn VGND VGND VPWR VPWR _14097_/A sky130_fd_sc_hd__dfrtp_4
X_22423_ _16345_/Y _22677_/B _22422_/X _16054_/Y _22265_/X VGND VGND VPWR VPWR _22423_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_109_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22295__B1 _22885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12783__B1 _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25142_ _24109_/CLK _14371_/X HRESETn VGND VGND VPWR VPWR _25142_/Q sky130_fd_sc_hd__dfrtp_4
X_22354_ _22055_/X _22354_/B VGND VGND VPWR VPWR _22354_/X sky130_fd_sc_hd__or2_4
XFILLER_136_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21305_ _17206_/X _21303_/X _13122_/A _21304_/X VGND VGND VPWR VPWR _21305_/X sky130_fd_sc_hd__a2bb2o_4
X_25073_ _25070_/CLK _25073_/D HRESETn VGND VGND VPWR VPWR _13573_/A sky130_fd_sc_hd__dfrtp_4
X_22285_ _21295_/X VGND VGND VPWR VPWR _22396_/C sky130_fd_sc_hd__buf_2
XANTENNA__22779__A1_N _12440_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24024_ _24055_/CLK _24024_/D HRESETn VGND VGND VPWR VPWR _13118_/A sky130_fd_sc_hd__dfrtp_4
X_21236_ _21253_/A _19102_/Y VGND VGND VPWR VPWR _21236_/X sky130_fd_sc_hd__or2_4
XFILLER_105_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16277__A1 _15669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21167_ _24199_/Q VGND VGND VPWR VPWR _21184_/A sky130_fd_sc_hd__buf_2
XFILLER_137_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17317__C _17253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20118_ _20105_/X VGND VGND VPWR VPWR _20118_/X sky130_fd_sc_hd__buf_2
XFILLER_131_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24352__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21098_ _21098_/A VGND VGND VPWR VPWR _21098_/X sky130_fd_sc_hd__buf_2
XFILLER_28_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12940_ _12761_/Y _12600_/X VGND VGND VPWR VPWR _12979_/B sky130_fd_sc_hd__or2_4
X_20049_ _23514_/Q VGND VGND VPWR VPWR _22068_/B sky130_fd_sc_hd__inv_2
X_24926_ _24926_/CLK _24926_/D HRESETn VGND VGND VPWR VPWR _11729_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_86_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12871_ _12871_/A _12871_/B VGND VGND VPWR VPWR _12873_/B sky130_fd_sc_hd__or2_4
X_24857_ _24865_/CLK _15744_/X HRESETn VGND VGND VPWR VPWR _24857_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20781__B1 _20706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14610_ _14610_/A _25070_/Q VGND VGND VPWR VPWR _14610_/X sky130_fd_sc_hd__or2_4
X_11822_ _11821_/X VGND VGND VPWR VPWR _11822_/X sky130_fd_sc_hd__buf_2
XFILLER_27_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23808_ _23832_/CLK _23808_/D VGND VGND VPWR VPWR _19208_/A sky130_fd_sc_hd__dfxtp_4
X_15590_ _24899_/Q VGND VGND VPWR VPWR _15590_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14460__B1 _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24788_ _24832_/CLK _15889_/X HRESETn VGND VGND VPWR VPWR _24788_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _11753_/A VGND VGND VPWR VPWR _11753_/Y sky130_fd_sc_hd__inv_2
X_14541_ _14541_/A _14540_/X VGND VGND VPWR VPWR _25088_/D sky130_fd_sc_hd__or2_4
XFILLER_81_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23739_ _23887_/CLK _19405_/X VGND VGND VPWR VPWR _23739_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17260_/A _17260_/B VGND VGND VPWR VPWR _17260_/X sky130_fd_sc_hd__or2_4
XPHY_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11682_/A _24214_/Q _11682_/Y _11683_/Y VGND VGND VPWR VPWR _11684_/X sky130_fd_sc_hd__o22a_4
X_14472_ _25109_/Q VGND VGND VPWR VPWR _14472_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23078__A2 _21287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _22992_/A VGND VGND VPWR VPWR _16211_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25140__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ _13455_/A _23630_/Q VGND VGND VPWR VPWR _13425_/B sky130_fd_sc_hd__or2_4
XANTENNA__13589__A _13588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22286__B1 _12514_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25409_ _25400_/CLK _25409_/D HRESETn VGND VGND VPWR VPWR _25409_/Q sky130_fd_sc_hd__dfrtp_4
X_17191_ _17183_/X _17191_/B _17187_/X _17191_/D VGND VGND VPWR VPWR _17202_/C sky130_fd_sc_hd__or4_4
XFILLER_128_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22825__A2 _22824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13354_ _13386_/A _13354_/B _13354_/C VGND VGND VPWR VPWR _13358_/B sky130_fd_sc_hd__and3_4
X_16142_ _22484_/A VGND VGND VPWR VPWR _16142_/Y sky130_fd_sc_hd__inv_2
X_12305_ _12305_/A VGND VGND VPWR VPWR _12305_/Y sky130_fd_sc_hd__inv_2
X_13285_ _13390_/A _13285_/B _13284_/X VGND VGND VPWR VPWR _13285_/X sky130_fd_sc_hd__or3_4
X_16073_ _24704_/Q VGND VGND VPWR VPWR _16073_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15712__B1 _24873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12236_ _12235_/X _24747_/Q _12235_/A _24747_/Q VGND VGND VPWR VPWR _12236_/X sky130_fd_sc_hd__a2bb2o_4
X_15024_ _25000_/Q _14991_/Y _25005_/Q _15023_/Y VGND VGND VPWR VPWR _15024_/X sky130_fd_sc_hd__a2bb2o_4
X_19901_ _19901_/A VGND VGND VPWR VPWR _21669_/B sky130_fd_sc_hd__inv_2
Xclkbuf_4_9_0_HCLK clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12940__B _12600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19832_ _19831_/Y _19829_/X _19787_/X _19829_/X VGND VGND VPWR VPWR _19832_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11837__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12167_ _12121_/A _14325_/A _12166_/X _12163_/A VGND VGND VPWR VPWR _12167_/X sky130_fd_sc_hd__a211o_4
XFILLER_69_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19763_ _13362_/B VGND VGND VPWR VPWR _19763_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24093__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12098_ _12097_/X VGND VGND VPWR VPWR _13496_/B sky130_fd_sc_hd__buf_2
X_16975_ _24711_/Q _24368_/Q _16054_/Y _17038_/B VGND VGND VPWR VPWR _16980_/B sky130_fd_sc_hd__o22a_4
X_18714_ _18738_/A _18714_/B _18713_/X VGND VGND VPWR VPWR _24142_/D sky130_fd_sc_hd__and3_4
X_15926_ _15655_/X _15835_/X _15845_/X _12983_/A _15925_/X VGND VGND VPWR VPWR _15926_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_77_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24022__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19694_ _23640_/Q VGND VGND VPWR VPWR _19694_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_5_30_0_HCLK clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18645_ _18638_/X _18642_/X _18643_/X _18645_/D VGND VGND VPWR VPWR _18645_/X sky130_fd_sc_hd__or4_4
XANTENNA__21046__A _21015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15857_ _15857_/A VGND VGND VPWR VPWR _15857_/X sky130_fd_sc_hd__buf_2
X_14808_ _14807_/X VGND VGND VPWR VPWR _14809_/A sky130_fd_sc_hd__buf_2
XANTENNA__25299__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18576_ _18555_/A _18576_/B _18575_/Y VGND VGND VPWR VPWR _24152_/D sky130_fd_sc_hd__and3_4
XFILLER_75_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15788_ _15795_/A VGND VGND VPWR VPWR _15788_/X sky130_fd_sc_hd__buf_2
XANTENNA__15794__A3 _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17527_ _17527_/A VGND VGND VPWR VPWR _17578_/C sky130_fd_sc_hd__inv_2
XANTENNA__25228__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14739_ _14731_/X _14738_/Y _25054_/Q _14723_/Y VGND VGND VPWR VPWR _14739_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19390__B1 _19389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17458_ _17456_/A _17457_/A _17456_/Y _17457_/Y VGND VGND VPWR VPWR _17458_/X sky130_fd_sc_hd__o22a_4
X_16409_ _15118_/Y _16406_/X _16408_/X _16406_/X VGND VGND VPWR VPWR _24585_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14754__A1 _21612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17389_ _17389_/A _17388_/X VGND VGND VPWR VPWR _20620_/B sky130_fd_sc_hd__or2_4
XANTENNA__15951__B1 _24758_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19142__B1 _19117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19128_ _19014_/A _19038_/B _19399_/C VGND VGND VPWR VPWR _19129_/A sky130_fd_sc_hd__or3_4
XFILLER_119_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_154_0_HCLK clkbuf_7_77_0_HCLK/X VGND VGND VPWR VPWR _24186_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22292__A3 _22287_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19059_ _19058_/Y _19052_/X _19010_/X _19052_/A VGND VGND VPWR VPWR _19059_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24863__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22070_ _14680_/X VGND VGND VPWR VPWR _22070_/X sky130_fd_sc_hd__buf_2
X_21021_ _22523_/A VGND VGND VPWR VPWR _21021_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17208__B1 _16352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22972_ _21111_/X VGND VGND VPWR VPWR _22972_/X sky130_fd_sc_hd__buf_2
XFILLER_110_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18956__B1 _18955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24711_ _24712_/CLK _16055_/X HRESETn VGND VGND VPWR VPWR _24711_/Q sky130_fd_sc_hd__dfrtp_4
X_21923_ _21944_/A _20347_/Y VGND VGND VPWR VPWR _21923_/X sky130_fd_sc_hd__or2_4
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21854_ _21098_/A _21854_/B _21854_/C VGND VGND VPWR VPWR _21862_/C sky130_fd_sc_hd__and3_4
X_24642_ _24643_/CLK _24642_/D HRESETn VGND VGND VPWR VPWR _16249_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_93_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21307__A2 _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20805_ _20803_/Y _20800_/X _20804_/X VGND VGND VPWR VPWR _20805_/X sky130_fd_sc_hd__o21a_4
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21785_ _21449_/A _19504_/Y VGND VGND VPWR VPWR _21785_/X sky130_fd_sc_hd__or2_4
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24573_ _24596_/CLK _24573_/D HRESETn VGND VGND VPWR VPWR _15077_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20736_ _20734_/Y _20731_/Y _20740_/B VGND VGND VPWR VPWR _20736_/X sky130_fd_sc_hd__o21a_4
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23524_ _23394_/CLK _20025_/X VGND VGND VPWR VPWR _23524_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_50_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23455_ _23478_/CLK _23455_/D VGND VGND VPWR VPWR _23455_/Q sky130_fd_sc_hd__dfxtp_4
X_20667_ _20488_/B VGND VGND VPWR VPWR _20667_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21122__C _14406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22406_ _16702_/Y _22406_/B VGND VGND VPWR VPWR _22406_/X sky130_fd_sc_hd__and2_4
XFILLER_104_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23386_ _24219_/CLK _20384_/X VGND VGND VPWR VPWR _23386_/Q sky130_fd_sc_hd__dfxtp_4
X_20598_ _20593_/X _20597_/X _14089_/X VGND VGND VPWR VPWR _20598_/X sky130_fd_sc_hd__o21a_4
XFILLER_109_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22515__A _21024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22337_ _21912_/X _22337_/B _22337_/C VGND VGND VPWR VPWR _22337_/X sky130_fd_sc_hd__and3_4
X_25125_ _25101_/CLK _25125_/D HRESETn VGND VGND VPWR VPWR _25125_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__17609__A _17885_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16513__A _24544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13070_ _13042_/A VGND VGND VPWR VPWR _13076_/A sky130_fd_sc_hd__buf_2
X_25056_ _25055_/CLK _25056_/D HRESETn VGND VGND VPWR VPWR _21643_/A sky130_fd_sc_hd__dfrtp_4
X_22268_ _22407_/B VGND VGND VPWR VPWR _22268_/X sky130_fd_sc_hd__buf_2
XANTENNA__24533__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12021_ _12021_/A VGND VGND VPWR VPWR _12021_/Y sky130_fd_sc_hd__inv_2
X_24007_ _24041_/CLK _20727_/X HRESETn VGND VGND VPWR VPWR _24007_/Q sky130_fd_sc_hd__dfrtp_4
X_21219_ _21112_/B _21216_/X _21323_/A _21218_/Y VGND VGND VPWR VPWR _21220_/C sky130_fd_sc_hd__a211o_4
XFILLER_65_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22199_ _21238_/X _22197_/X _22198_/X VGND VGND VPWR VPWR _22199_/X sky130_fd_sc_hd__and3_4
XFILLER_116_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16760_ _15003_/Y _16759_/X _15739_/X _16759_/X VGND VGND VPWR VPWR _16760_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13972_ scl_oen_o_S5 _13966_/X _13967_/Y _13971_/Y VGND VGND VPWR VPWR _13973_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_76_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22743__A1 _21280_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15711_ _15711_/A VGND VGND VPWR VPWR _15711_/X sky130_fd_sc_hd__buf_2
X_12923_ _12922_/X VGND VGND VPWR VPWR _25371_/D sky130_fd_sc_hd__inv_2
X_24909_ _24909_/CLK _24909_/D HRESETn VGND VGND VPWR VPWR _15565_/A sky130_fd_sc_hd__dfrtp_4
X_16691_ _22634_/A _16688_/X _15750_/X _16688_/X VGND VGND VPWR VPWR _24478_/D sky130_fd_sc_hd__a2bb2o_4
X_18430_ _16230_/Y _24159_/Q _16230_/Y _24159_/Q VGND VGND VPWR VPWR _18431_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25392__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15642_ _15642_/A _22824_/A VGND VGND VPWR VPWR _16640_/B sky130_fd_sc_hd__or2_4
X_12854_ _12854_/A _12854_/B VGND VGND VPWR VPWR _12877_/B sky130_fd_sc_hd__or2_4
XANTENNA__25321__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11805_ _11794_/X VGND VGND VPWR VPWR _11805_/X sky130_fd_sc_hd__buf_2
X_18361_ _18361_/A VGND VGND VPWR VPWR _18361_/Y sky130_fd_sc_hd__inv_2
X_15573_ _15572_/Y _15568_/X _11761_/X _15568_/X VGND VGND VPWR VPWR _15573_/X sky130_fd_sc_hd__a2bb2o_4
X_12785_ _24781_/Q VGND VGND VPWR VPWR _12785_/Y sky130_fd_sc_hd__inv_2
XPHY_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17177_/A _17311_/Y VGND VGND VPWR VPWR _17312_/X sky130_fd_sc_hd__or2_4
XFILLER_30_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14524_ _21841_/A _14511_/X _21709_/A _14513_/X VGND VGND VPWR VPWR _14524_/X sky130_fd_sc_hd__o22a_4
XFILLER_42_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11736_ _21018_/A VGND VGND VPWR VPWR _21582_/B sky130_fd_sc_hd__buf_2
X_18292_ _21192_/A VGND VGND VPWR VPWR _18293_/B sky130_fd_sc_hd__buf_2
XPHY_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _17240_/Y _17365_/A _17348_/A _17243_/D VGND VGND VPWR VPWR _17243_/X sky130_fd_sc_hd__or4_4
XFILLER_109_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ _14452_/X _14454_/X _14411_/X _14454_/X VGND VGND VPWR VPWR _14455_/X sky130_fd_sc_hd__a2bb2o_4
X_11667_ _11667_/A VGND VGND VPWR VPWR _13718_/A sky130_fd_sc_hd__inv_2
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _13301_/X _13404_/X _13405_/X VGND VGND VPWR VPWR _13406_/X sky130_fd_sc_hd__and3_4
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17174_ _17174_/A VGND VGND VPWR VPWR _17246_/C sky130_fd_sc_hd__inv_2
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14386_ _14386_/A VGND VGND VPWR VPWR _14386_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22274__A3 _21290_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12211__A2 _22400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22425__A _22425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_227_0_HCLK clkbuf_8_227_0_HCLK/A VGND VGND VPWR VPWR _24800_/CLK sky130_fd_sc_hd__clkbuf_1
X_16125_ _16087_/A VGND VGND VPWR VPWR _16125_/X sky130_fd_sc_hd__buf_2
X_13337_ _17452_/B _13337_/B VGND VGND VPWR VPWR _13337_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_4_7_0_HCLK_A clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22144__B _22654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16056_ _24710_/Q VGND VGND VPWR VPWR _16056_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24274__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13268_ _13454_/A _13264_/X _13267_/X VGND VGND VPWR VPWR _13268_/X sky130_fd_sc_hd__or3_4
X_15007_ _15063_/B VGND VGND VPWR VPWR _15251_/B sky130_fd_sc_hd__buf_2
X_12219_ _25429_/Q VGND VGND VPWR VPWR _12220_/A sky130_fd_sc_hd__inv_2
XANTENNA__22431__B1 _12536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24203__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13199_ _11964_/X VGND VGND VPWR VPWR _13199_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19815_ _19802_/Y VGND VGND VPWR VPWR _19815_/X sky130_fd_sc_hd__buf_2
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17254__A _17254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16958_ _16046_/Y _24371_/Q _16046_/Y _24371_/Q VGND VGND VPWR VPWR _16958_/X sky130_fd_sc_hd__a2bb2o_4
X_19746_ _19745_/Y _19743_/X _19700_/X _19743_/X VGND VGND VPWR VPWR _19746_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18938__B1 _16852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15909_ _12795_/Y _15904_/X _15840_/X _15868_/X VGND VGND VPWR VPWR _15909_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25409__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19677_ _19675_/Y _19676_/X _19553_/X _19676_/X VGND VGND VPWR VPWR _23647_/D sky130_fd_sc_hd__a2bb2o_4
X_16889_ _16887_/Y _16880_/X _16888_/X _16880_/A VGND VGND VPWR VPWR _16889_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18628_ _24142_/Q VGND VGND VPWR VPWR _18705_/A sky130_fd_sc_hd__inv_2
XFILLER_25_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15767__A3 _15766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21504__A _21504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25062__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18559_ _18472_/A _18418_/Y _18475_/C _18592_/A VGND VGND VPWR VPWR _18559_/X sky130_fd_sc_hd__or4_4
X_21570_ _22123_/A VGND VGND VPWR VPWR _21570_/X sky130_fd_sc_hd__buf_2
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_37_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_75_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20521_ _24069_/Q _20519_/X _20493_/X VGND VGND VPWR VPWR _20521_/X sky130_fd_sc_hd__a21o_4
XFILLER_53_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19115__B1 _19071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23240_ _23208_/A _23231_/Y _23235_/X _23240_/D VGND VGND VPWR VPWR _23240_/X sky130_fd_sc_hd__or4_4
X_20452_ _20452_/A _20452_/B VGND VGND VPWR VPWR _20452_/X sky130_fd_sc_hd__and2_4
XFILLER_88_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23171_ _24593_/Q _23171_/B VGND VGND VPWR VPWR _23175_/B sky130_fd_sc_hd__or2_4
X_20383_ _18237_/A VGND VGND VPWR VPWR _20383_/X sky130_fd_sc_hd__buf_2
XFILLER_107_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22122_ _21529_/X _22121_/X _21532_/X _24847_/Q _21533_/X VGND VGND VPWR VPWR _22122_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_133_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22053_ _21890_/X _22053_/B _22052_/X VGND VGND VPWR VPWR _22053_/X sky130_fd_sc_hd__and3_4
XFILLER_115_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21004_ _21053_/A _21004_/B VGND VGND VPWR VPWR _21004_/X sky130_fd_sc_hd__and2_4
XFILLER_134_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12910__B1 _12874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23166__A _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23997__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23926__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22955_ _22714_/X _22955_/B VGND VGND VPWR VPWR _22955_/Y sky130_fd_sc_hd__nor2_4
XFILLER_16_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21906_ _21886_/A _21906_/B VGND VGND VPWR VPWR _21906_/X sky130_fd_sc_hd__or2_4
XFILLER_16_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14415__B1 _14414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_119_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_239_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22886_ _24451_/Q _22421_/X _22885_/X VGND VGND VPWR VPWR _22886_/X sky130_fd_sc_hd__o21a_4
XFILLER_55_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24625_ _24355_/CLK _24625_/D HRESETn VGND VGND VPWR VPWR _16295_/A sky130_fd_sc_hd__dfrtp_4
X_21837_ _21837_/A _22695_/B _22695_/C VGND VGND VPWR VPWR _21837_/X sky130_fd_sc_hd__and3_4
XANTENNA__19505__A2_N _19500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12570_ _12570_/A VGND VGND VPWR VPWR _12570_/Y sky130_fd_sc_hd__inv_2
X_21768_ _21763_/X _21766_/X _21767_/X VGND VGND VPWR VPWR _21768_/X sky130_fd_sc_hd__o21a_4
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24556_ _24557_/CLK _16484_/X HRESETn VGND VGND VPWR VPWR _24556_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20719_ _22513_/A _20698_/X _20706_/X _20718_/X VGND VGND VPWR VPWR _20719_/X sky130_fd_sc_hd__o22a_4
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23507_ _24208_/CLK _20068_/X VGND VGND VPWR VPWR _23507_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24785__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21699_ _21699_/A VGND VGND VPWR VPWR _21699_/Y sky130_fd_sc_hd__inv_2
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24487_ _24487_/CLK _24487_/D HRESETn VGND VGND VPWR VPWR _24487_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240_ _14238_/Y _14236_/X _14239_/X _14236_/X VGND VGND VPWR VPWR _14240_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24714__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23438_ _23904_/CLK _23438_/D VGND VGND VPWR VPWR _23438_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14171_ _25197_/Q _23950_/Q VGND VGND VPWR VPWR _14171_/X sky130_fd_sc_hd__or2_4
XANTENNA__22661__B1 _17759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23369_ _24496_/CLK _20812_/A VGND VGND VPWR VPWR _13670_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_5_0_0_HCLK_A clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13122_ _13122_/A _23997_/Q VGND VGND VPWR VPWR _13123_/B sky130_fd_sc_hd__nor2_4
X_25108_ _24945_/CLK _25108_/D HRESETn VGND VGND VPWR VPWR _14474_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_106_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23205__A2 _22998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_57_0_HCLK clkbuf_8_57_0_HCLK/A VGND VGND VPWR VPWR _25255_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_79_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13053_ _12358_/Y _13052_/X VGND VGND VPWR VPWR _13067_/B sky130_fd_sc_hd__or2_4
X_17930_ _17930_/A _23868_/Q VGND VGND VPWR VPWR _17931_/C sky130_fd_sc_hd__or2_4
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25039_ _24070_/CLK _14840_/X HRESETn VGND VGND VPWR VPWR _25039_/Q sky130_fd_sc_hd__dfrtp_4
X_12004_ _11992_/X VGND VGND VPWR VPWR _12004_/Y sky130_fd_sc_hd__inv_2
X_17861_ _16918_/A _17861_/B VGND VGND VPWR VPWR _17863_/B sky130_fd_sc_hd__or2_4
XFILLER_132_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18632__A2 _18630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16812_ _14919_/Y _16807_/X HWDATA[24] _16811_/X VGND VGND VPWR VPWR _24425_/D sky130_fd_sc_hd__a2bb2o_4
X_19600_ _19598_/Y _19593_/X _19599_/X _19593_/X VGND VGND VPWR VPWR _23672_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17792_ _16943_/Y _17792_/B _17792_/C VGND VGND VPWR VPWR _17792_/X sky130_fd_sc_hd__or3_4
X_19531_ _19530_/Y _19528_/X _11955_/X _19528_/X VGND VGND VPWR VPWR _19531_/X sky130_fd_sc_hd__a2bb2o_4
X_16743_ _16739_/A VGND VGND VPWR VPWR _16743_/X sky130_fd_sc_hd__buf_2
XANTENNA__25502__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13955_ _13921_/Y _13930_/D _13947_/A VGND VGND VPWR VPWR _13960_/A sky130_fd_sc_hd__or3_4
XFILLER_46_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15306__B _15336_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12906_ _12905_/X VGND VGND VPWR VPWR _12906_/Y sky130_fd_sc_hd__inv_2
X_19462_ _19055_/X VGND VGND VPWR VPWR _19462_/X sky130_fd_sc_hd__buf_2
XFILLER_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16674_ _16673_/Y _16671_/X _16405_/X _16671_/X VGND VGND VPWR VPWR _24485_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13886_ _23987_/Q VGND VGND VPWR VPWR _13886_/X sky130_fd_sc_hd__buf_2
XFILLER_35_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18413_ _18413_/A _18408_/X _18413_/C _18412_/X VGND VGND VPWR VPWR _18413_/X sky130_fd_sc_hd__or4_4
X_15625_ _15625_/A VGND VGND VPWR VPWR _15625_/Y sky130_fd_sc_hd__inv_2
X_12837_ _12791_/X _12836_/X VGND VGND VPWR VPWR _12838_/A sky130_fd_sc_hd__or2_4
X_19393_ _19391_/Y _19392_/X _19370_/X _19392_/X VGND VGND VPWR VPWR _19393_/X sky130_fd_sc_hd__a2bb2o_4
X_18344_ _18344_/A _18338_/X VGND VGND VPWR VPWR _18344_/X sky130_fd_sc_hd__and2_4
X_15556_ _22695_/B VGND VGND VPWR VPWR _16640_/A sky130_fd_sc_hd__buf_2
X_12768_ _12846_/B VGND VGND VPWR VPWR _12944_/B sky130_fd_sc_hd__buf_2
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14507_ _14505_/X _14517_/A _20441_/B VGND VGND VPWR VPWR _14507_/X sky130_fd_sc_hd__a21o_4
XANTENNA__14709__A1 _21781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11719_ _15991_/A _11719_/B _15991_/C _15991_/D VGND VGND VPWR VPWR _11720_/B sky130_fd_sc_hd__or4_4
X_18275_ _18275_/A VGND VGND VPWR VPWR _18275_/X sky130_fd_sc_hd__buf_2
XFILLER_124_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15906__B1 _24776_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15487_ _24063_/D _15486_/X VGND VGND VPWR VPWR _15487_/X sky130_fd_sc_hd__or2_4
X_12699_ _12565_/Y _12693_/X _12695_/Y _12653_/X VGND VGND VPWR VPWR _12699_/X sky130_fd_sc_hd__a211o_4
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17226_ _16284_/Y _24358_/Q _16284_/Y _24358_/Q VGND VGND VPWR VPWR _17229_/B sky130_fd_sc_hd__a2bb2o_4
X_14438_ _22302_/A _14437_/X _14411_/X _14437_/X VGND VGND VPWR VPWR _25124_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24455__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13777__A _13777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17157_ _17156_/A _17160_/A VGND VGND VPWR VPWR _17157_/X sky130_fd_sc_hd__or2_4
XANTENNA__22652__B1 _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14369_ _14354_/Y _14368_/X _25468_/Q _14360_/X VGND VGND VPWR VPWR _25143_/D sky130_fd_sc_hd__o22a_4
XFILLER_7_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16108_ _23043_/A VGND VGND VPWR VPWR _16108_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13496__B _13496_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17088_ _17384_/B _17088_/B _17087_/X VGND VGND VPWR VPWR _17089_/A sky130_fd_sc_hd__or3_4
XANTENNA__16331__B1 _16231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16039_ _24717_/Q VGND VGND VPWR VPWR _16039_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15992__A _16371_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22404__B1 _22270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25243__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19729_ _19729_/A VGND VGND VPWR VPWR _19729_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22740_ _24750_/Q _22626_/B VGND VGND VPWR VPWR _22740_/X sky130_fd_sc_hd__or2_4
XFILLER_25_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22671_ _22671_/A _22671_/B VGND VGND VPWR VPWR _22671_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__14948__B2 _24413_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12856__A _12602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11760__A _11777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21622_ _21622_/A VGND VGND VPWR VPWR _21623_/A sky130_fd_sc_hd__buf_2
X_24410_ _24998_/CLK _16841_/X HRESETn VGND VGND VPWR VPWR _14934_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25390_ _25411_/CLK _12734_/X HRESETn VGND VGND VPWR VPWR _25390_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21553_ _14209_/Y _14194_/A _14235_/Y _14221_/A VGND VGND VPWR VPWR _21554_/A sky130_fd_sc_hd__o22a_4
XFILLER_21_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24341_ _24355_/CLK _24341_/D HRESETn VGND VGND VPWR VPWR _17248_/A sky130_fd_sc_hd__dfrtp_4
X_20504_ _20490_/A _20504_/B _20504_/C VGND VGND VPWR VPWR _20504_/X sky130_fd_sc_hd__or3_4
XANTENNA__24076__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24272_ _24267_/CLK _24272_/D HRESETn VGND VGND VPWR VPWR _17785_/A sky130_fd_sc_hd__dfrtp_4
X_21484_ _21484_/A _19530_/Y VGND VGND VPWR VPWR _21484_/X sky130_fd_sc_hd__or2_4
XANTENNA__24196__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23223_ _12385_/B _21524_/X _24273_/Q _22483_/X VGND VGND VPWR VPWR _23223_/X sky130_fd_sc_hd__a2bb2o_4
X_20435_ _20444_/A _20433_/X VGND VGND VPWR VPWR _20437_/C sky130_fd_sc_hd__and2_4
XFILLER_10_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17495__A1_N _25513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24125__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16063__A _24708_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_210_0_HCLK clkbuf_8_211_0_HCLK/A VGND VGND VPWR VPWR _24492_/CLK sky130_fd_sc_hd__clkbuf_1
X_23154_ _23105_/X _23149_/Y _23150_/X _23153_/X VGND VGND VPWR VPWR _23154_/X sky130_fd_sc_hd__a2bb2o_4
X_20366_ _20360_/Y VGND VGND VPWR VPWR _20366_/X sky130_fd_sc_hd__buf_2
XFILLER_101_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22105_ _22102_/X _22104_/X _21306_/A VGND VGND VPWR VPWR _22105_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_136_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15676__A2 _15669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23085_ _23085_/A _23082_/X _23085_/C VGND VGND VPWR VPWR _23085_/X sky130_fd_sc_hd__and3_4
X_20297_ _18275_/A _19971_/X _20276_/C VGND VGND VPWR VPWR _20298_/A sky130_fd_sc_hd__or3_4
XANTENNA__22512__B _21428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22036_ _22036_/A _19604_/Y VGND VGND VPWR VPWR _22036_/X sky130_fd_sc_hd__and2_4
XANTENNA__22946__B2 _22827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21409__A _21409_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11935__A _11947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23987_ _24070_/CLK _23987_/D HRESETn VGND VGND VPWR VPWR _23987_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13740_ _13740_/A VGND VGND VPWR VPWR _13743_/A sky130_fd_sc_hd__inv_2
XANTENNA__17622__A _17885_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22938_ _22808_/X _22935_/X _22938_/C VGND VGND VPWR VPWR _22938_/X sky130_fd_sc_hd__and3_4
XFILLER_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13671_ _24877_/Q VGND VGND VPWR VPWR _13671_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24966__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22869_ _12199_/Y _22489_/X _24263_/Q _21045_/X VGND VGND VPWR VPWR _22869_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16238__A _11812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15410_ _24968_/Q _15409_/Y VGND VGND VPWR VPWR _15411_/B sky130_fd_sc_hd__or2_4
X_12622_ _12622_/A _12645_/A _12636_/A _12642_/B VGND VGND VPWR VPWR _12623_/C sky130_fd_sc_hd__or4_4
XFILLER_58_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24608_ _24177_/CLK _24608_/D HRESETn VGND VGND VPWR VPWR _22478_/A sky130_fd_sc_hd__dfrtp_4
X_16390_ _16388_/Y _16389_/X _16297_/X _16389_/X VGND VGND VPWR VPWR _16390_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21134__B1 _23344_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15341_ _15080_/Y _15338_/X _15340_/Y VGND VGND VPWR VPWR _24988_/D sky130_fd_sc_hd__o21a_4
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ _25390_/Q _12552_/A _12729_/A _12552_/Y VGND VGND VPWR VPWR _12557_/C sky130_fd_sc_hd__o22a_4
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24539_ _24541_/CLK _16529_/X HRESETn VGND VGND VPWR VPWR _24539_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18060_ _15695_/X _18040_/X _18059_/X _24235_/Q _18019_/X VGND VGND VPWR VPWR _18060_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_20_0_HCLK clkbuf_6_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_41_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15272_ _15272_/A VGND VGND VPWR VPWR _15272_/Y sky130_fd_sc_hd__inv_2
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ _12503_/A _12482_/X _12483_/X VGND VGND VPWR VPWR _25429_/D sky130_fd_sc_hd__and3_4
XANTENNA__16561__B1 _16300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17011_ _17004_/X _17011_/B _17008_/X _17010_/X VGND VGND VPWR VPWR _17017_/C sky130_fd_sc_hd__or4_4
XANTENNA__12178__B2 _24746_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14223_ _14223_/A _14223_/B VGND VGND VPWR VPWR _14224_/A sky130_fd_sc_hd__nor2_4
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18302__A1 _18299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14154_ _14154_/A VGND VGND VPWR VPWR _14154_/Y sky130_fd_sc_hd__inv_2
X_13105_ _13105_/A VGND VGND VPWR VPWR _13105_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14085_ _13982_/A _14081_/X _14078_/X _13980_/A _14084_/X VGND VGND VPWR VPWR _14085_/X
+ sky130_fd_sc_hd__a32o_4
X_18962_ _18959_/Y _18960_/X _18961_/X _18960_/X VGND VGND VPWR VPWR _23895_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22937__A1 _24522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13036_ _13029_/B VGND VGND VPWR VPWR _13037_/B sky130_fd_sc_hd__inv_2
X_17913_ _15684_/A _14769_/X _15915_/X _17912_/X VGND VGND VPWR VPWR _17920_/C sky130_fd_sc_hd__a211o_4
XFILLER_117_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18893_ _23995_/Q _14535_/Y _20982_/A _20531_/A VGND VGND VPWR VPWR _24105_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22401__A3 _22130_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12350__B2 _24821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11845__A HWDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17844_ _17844_/A VGND VGND VPWR VPWR _17844_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17775_ _16948_/X _17765_/D VGND VGND VPWR VPWR _17776_/A sky130_fd_sc_hd__or2_4
X_14987_ _15199_/A VGND VGND VPWR VPWR _15190_/A sky130_fd_sc_hd__buf_2
XANTENNA__18628__A _24142_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16726_ _15310_/B _16725_/X _16720_/X _16725_/X VGND VGND VPWR VPWR _24465_/D sky130_fd_sc_hd__a2bb2o_4
X_19514_ _20000_/C _18287_/X _18275_/A _18280_/X VGND VGND VPWR VPWR _19515_/A sky130_fd_sc_hd__or4_4
X_13938_ _13952_/A _13957_/B VGND VGND VPWR VPWR _13939_/B sky130_fd_sc_hd__nand2_4
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16919__A2 _16918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19445_ _14656_/Y _19152_/D _19013_/X VGND VGND VPWR VPWR _19445_/X sky130_fd_sc_hd__or3_4
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16657_ _24491_/Q VGND VGND VPWR VPWR _23120_/A sky130_fd_sc_hd__inv_2
X_13869_ _22172_/A _13861_/X _22111_/A _13863_/X VGND VGND VPWR VPWR _13869_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_102_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_205_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15608_ _15607_/Y _15605_/X _11813_/X _15605_/X VGND VGND VPWR VPWR _15608_/X sky130_fd_sc_hd__a2bb2o_4
X_19376_ _17946_/B VGND VGND VPWR VPWR _19376_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16588_ _16583_/A VGND VGND VPWR VPWR _16588_/X sky130_fd_sc_hd__buf_2
XANTENNA__24636__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18327_ _24197_/Q VGND VGND VPWR VPWR _19728_/A sky130_fd_sc_hd__buf_2
X_15539_ _13789_/D _15535_/X HADDR[2] _15538_/X VGND VGND VPWR VPWR _24914_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14891__A _25022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18258_ _18235_/A _18253_/X _16270_/X _24213_/Q _18231_/A VGND VGND VPWR VPWR _24213_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_72_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16552__B1 _16380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12169__A1 _12123_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17209_ _16334_/Y _24340_/Q _16334_/Y _24340_/Q VGND VGND VPWR VPWR _17211_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18189_ _18054_/X _18189_/B VGND VGND VPWR VPWR _18189_/X sky130_fd_sc_hd__or2_4
X_20220_ _20219_/Y _20217_/X _19715_/X _20217_/X VGND VGND VPWR VPWR _23449_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16304__B1 _15949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11739__B _22913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20151_ _23475_/Q VGND VGND VPWR VPWR _22197_/B sky130_fd_sc_hd__inv_2
XANTENNA__25495__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16611__A _16611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_40_0_HCLK clkbuf_7_20_0_HCLK/X VGND VGND VPWR VPWR _23828_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25424__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20082_ _16861_/A VGND VGND VPWR VPWR _20082_/X sky130_fd_sc_hd__buf_2
XANTENNA__20133__A _20140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23910_ _23478_/CLK _18917_/X VGND VGND VPWR VPWR _18916_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24890_ _24893_/CLK _15613_/X HRESETn VGND VGND VPWR VPWR _15611_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24940__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17280__A1 _17261_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23841_ _23854_/CLK _23841_/D VGND VGND VPWR VPWR _23841_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22156__A2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17442__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20984_ _20984_/A _23917_/Q VGND VGND VPWR VPWR _20984_/X sky130_fd_sc_hd__and2_4
X_23772_ _23772_/CLK _19314_/X VGND VGND VPWR VPWR _19309_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25511_ _25514_/CLK _11849_/X HRESETn VGND VGND VPWR VPWR _25511_/Q sky130_fd_sc_hd__dfrtp_4
X_22723_ _24448_/Q _22525_/X _22526_/X VGND VGND VPWR VPWR _22723_/X sky130_fd_sc_hd__o21a_4
XFILLER_80_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25442_ _25449_/CLK _25442_/D HRESETn VGND VGND VPWR VPWR _12252_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24377__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22654_ _22654_/A VGND VGND VPWR VPWR _22654_/X sky130_fd_sc_hd__buf_2
XANTENNA__16791__B1 _16717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21605_ _21609_/A _21605_/B _21605_/C VGND VGND VPWR VPWR _21605_/X sky130_fd_sc_hd__and3_4
XANTENNA__15897__A _11821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24306__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25373_ _24792_/CLK _12918_/X HRESETn VGND VGND VPWR VPWR _25373_/Q sky130_fd_sc_hd__dfrtp_4
X_22585_ _16594_/A _23226_/B _21731_/X _22584_/X VGND VGND VPWR VPWR _22586_/C sky130_fd_sc_hd__a211o_4
XFILLER_107_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22507__B _22613_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24324_ _23964_/CLK _17408_/X HRESETn VGND VGND VPWR VPWR _24324_/Q sky130_fd_sc_hd__dfstp_4
X_21536_ _12499_/A _22489_/A _24247_/Q _21422_/X VGND VGND VPWR VPWR _21536_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21467_ _21467_/A _21467_/B _21467_/C VGND VGND VPWR VPWR _21467_/X sky130_fd_sc_hd__and3_4
XANTENNA__20890__A2 _20884_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24255_ _24673_/CLK _24255_/D HRESETn VGND VGND VPWR VPWR _24255_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13210__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20418_ _15486_/X VGND VGND VPWR VPWR _20419_/B sky130_fd_sc_hd__inv_2
XANTENNA__22092__A1 _16611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23206_ _14905_/A _22135_/X _22997_/X _23205_/X VGND VGND VPWR VPWR _23207_/C sky130_fd_sc_hd__a211o_4
X_21398_ _21398_/A _21396_/X _21397_/X VGND VGND VPWR VPWR _21398_/X sky130_fd_sc_hd__and3_4
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18835__A2 _24142_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24186_ _24186_/CLK _18368_/X HRESETn VGND VGND VPWR VPWR _18365_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_135_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22523__A _22523_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20349_ _23399_/Q VGND VGND VPWR VPWR _21792_/B sky130_fd_sc_hd__inv_2
XFILLER_108_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23137_ _23065_/A _23137_/B _23136_/X VGND VGND VPWR VPWR _23138_/D sky130_fd_sc_hd__and3_4
XFILLER_122_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16521__A _16057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23941__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22919__A1 _13119_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22919__B2 _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23041__B1 _24726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23068_ _23068_/A _22722_/B VGND VGND VPWR VPWR _23071_/B sky130_fd_sc_hd__or2_4
XANTENNA__17336__B _17247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14910_ _14910_/A _14910_/B _14910_/C _14909_/X VGND VGND VPWR VPWR _14940_/B sky130_fd_sc_hd__or4_4
X_22019_ _22015_/X _22018_/X _21679_/X VGND VGND VPWR VPWR _22019_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_27_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15890_ _15886_/X _15887_/X _11800_/A _24787_/Q _15888_/X VGND VGND VPWR VPWR _24787_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_114_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16456__A2_N _16455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14841_ _14802_/A _14802_/B _14802_/A _14802_/B VGND VGND VPWR VPWR _14841_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23354__A _23338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19548__B1 _19547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17560_ _24304_/Q VGND VGND VPWR VPWR _17560_/Y sky130_fd_sc_hd__inv_2
X_14772_ _14772_/A _14772_/B _14769_/X _14771_/X VGND VGND VPWR VPWR _14772_/X sky130_fd_sc_hd__or4_4
XANTENNA__23073__B _22810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11984_ _11972_/X VGND VGND VPWR VPWR _11984_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16511_ _16504_/A VGND VGND VPWR VPWR _16511_/X sky130_fd_sc_hd__buf_2
X_13723_ _13685_/A _13685_/B VGND VGND VPWR VPWR _13723_/Y sky130_fd_sc_hd__nand2_4
X_17491_ _17491_/A VGND VGND VPWR VPWR _24310_/D sky130_fd_sc_hd__inv_2
XFILLER_72_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11843__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19230_ _19229_/Y _19227_/X _19206_/X _19227_/X VGND VGND VPWR VPWR _23801_/D sky130_fd_sc_hd__a2bb2o_4
X_16442_ _16442_/A VGND VGND VPWR VPWR _16442_/X sky130_fd_sc_hd__buf_2
XFILLER_32_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13654_ _13654_/A VGND VGND VPWR VPWR _13655_/B sky130_fd_sc_hd__inv_2
XFILLER_95_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12605_ _12665_/A VGND VGND VPWR VPWR _12693_/A sky130_fd_sc_hd__buf_2
X_19161_ _19159_/Y _19154_/X _19136_/X _19160_/X VGND VGND VPWR VPWR _23826_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16373_ _16373_/A _16728_/B VGND VGND VPWR VPWR _16381_/A sky130_fd_sc_hd__nor2_4
XANTENNA__22855__B1 _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24047__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _13846_/A _14560_/A _25242_/Q _14560_/B VGND VGND VPWR VPWR _13585_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18112_ _18176_/A _18112_/B _18112_/C VGND VGND VPWR VPWR _18113_/C sky130_fd_sc_hd__and3_4
XANTENNA__22417__B _22399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15324_ _15346_/A _15322_/X _15323_/X VGND VGND VPWR VPWR _24992_/D sky130_fd_sc_hd__and3_4
XANTENNA__15600__A _15588_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12536_ _24850_/Q VGND VGND VPWR VPWR _12536_/Y sky130_fd_sc_hd__inv_2
X_19092_ _22060_/B _19086_/X _16872_/X _19091_/X VGND VGND VPWR VPWR _19092_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16534__B1 _16359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18043_ _17999_/A _19044_/A VGND VGND VPWR VPWR _18044_/C sky130_fd_sc_hd__or2_4
X_15255_ _15282_/A _15253_/X _15254_/X VGND VGND VPWR VPWR _25006_/D sky130_fd_sc_hd__and3_4
X_12467_ _12509_/A VGND VGND VPWR VPWR _12503_/A sky130_fd_sc_hd__buf_2
XANTENNA__14216__A _20664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14206_ _14205_/Y _14199_/X _13840_/X _14201_/X VGND VGND VPWR VPWR _14206_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22083__A1 _21260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15186_ _25022_/Q _15185_/Y VGND VGND VPWR VPWR _15186_/X sky130_fd_sc_hd__or2_4
XANTENNA__22083__B2 _22082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12398_ _12398_/A VGND VGND VPWR VPWR _12398_/Y sky130_fd_sc_hd__inv_2
X_14137_ _14110_/X _14135_/X _25129_/Q _14136_/X VGND VGND VPWR VPWR _14137_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_113_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12571__B2 _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21830__B2 _17416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19994_ _23534_/Q VGND VGND VPWR VPWR _21479_/B sky130_fd_sc_hd__inv_2
Xclkbuf_7_27_0_HCLK clkbuf_7_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21049__A _22913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23032__B1 _24830_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14068_ _14007_/X _14065_/X _14057_/X _14001_/D _14066_/X VGND VGND VPWR VPWR _14068_/X
+ sky130_fd_sc_hd__a32o_4
X_18945_ _18333_/X _18335_/X _20231_/C _17462_/Y VGND VGND VPWR VPWR _18945_/X sky130_fd_sc_hd__or4_4
X_13019_ _13019_/A VGND VGND VPWR VPWR _25350_/D sky130_fd_sc_hd__inv_2
XFILLER_95_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18876_ _20566_/A _20566_/B VGND VGND VPWR VPWR _18876_/X sky130_fd_sc_hd__or2_4
XFILLER_94_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23927__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17827_ _17834_/A _17822_/X _17827_/C VGND VGND VPWR VPWR _17827_/X sky130_fd_sc_hd__and3_4
XANTENNA__12295__A1_N _12294_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24888__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16596__A1_N _16594_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13790__A _14406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12087__B1 _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17758_ _17758_/A _17758_/B _16914_/Y _17758_/D VGND VGND VPWR VPWR _17758_/X sky130_fd_sc_hd__or4_4
XANTENNA__24817__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16709_ _24470_/Q VGND VGND VPWR VPWR _16709_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11834__B1 _11833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17689_ _17662_/B _17688_/X VGND VGND VPWR VPWR _17689_/X sky130_fd_sc_hd__or2_4
XFILLER_90_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19428_ _17985_/B VGND VGND VPWR VPWR _19428_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24470__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21512__A _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19359_ _19358_/Y _19356_/X _19291_/X _19356_/X VGND VGND VPWR VPWR _23755_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16606__A _24509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22370_ _21616_/A _22370_/B VGND VGND VPWR VPWR _22370_/X sky130_fd_sc_hd__or2_4
XANTENNA__20128__A _20140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16534__A1_N _16533_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12853__B _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21321_ _15671_/A VGND VGND VPWR VPWR _22298_/B sky130_fd_sc_hd__buf_2
XFILLER_129_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21252_ _21252_/A _21252_/B VGND VGND VPWR VPWR _21254_/B sky130_fd_sc_hd__or2_4
XFILLER_89_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24040_ _24041_/CLK _24040_/D HRESETn VGND VGND VPWR VPWR _24040_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20203_ _20203_/A VGND VGND VPWR VPWR _20203_/X sky130_fd_sc_hd__buf_2
XFILLER_117_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21183_ _24200_/Q _21181_/X _21182_/X VGND VGND VPWR VPWR _21183_/X sky130_fd_sc_hd__and3_4
XFILLER_137_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20134_ _22071_/B _20128_/X _20085_/X _20133_/X VGND VGND VPWR VPWR _20134_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23023__B1 _12368_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19778__B1 _19777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20065_ _20065_/A _18325_/A VGND VGND VPWR VPWR _20065_/Y sky130_fd_sc_hd__nand2_4
XFILLER_57_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24942_ _24942_/CLK _15472_/X HRESETn VGND VGND VPWR VPWR _15470_/A sky130_fd_sc_hd__dfstp_4
XFILLER_135_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21585__B1 _22280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24873_ _24018_/CLK _15712_/X HRESETn VGND VGND VPWR VPWR _24873_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15264__B1 _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23824_ _25264_/CLK _23824_/D VGND VGND VPWR VPWR _18123_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24558__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23755_ _25503_/CLK _23755_/D VGND VGND VPWR VPWR _17967_/B sky130_fd_sc_hd__dfxtp_4
X_20967_ _20496_/C _22097_/A _14541_/A VGND VGND VPWR VPWR _20967_/X sky130_fd_sc_hd__a21o_4
XFILLER_109_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22706_ _22706_/A _21220_/A VGND VGND VPWR VPWR _22706_/X sky130_fd_sc_hd__or2_4
X_23686_ _23689_/CLK _23686_/D VGND VGND VPWR VPWR _19555_/A sky130_fd_sc_hd__dfxtp_4
X_20898_ _20896_/Y _20893_/X _20897_/X VGND VGND VPWR VPWR _20898_/X sky130_fd_sc_hd__o21a_4
XFILLER_41_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25425_ _25425_/CLK _25425_/D HRESETn VGND VGND VPWR VPWR _25425_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22837__B1 _22834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24140__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22637_ _22146_/A _22632_/X _21826_/X _22636_/Y VGND VGND VPWR VPWR _22638_/A sky130_fd_sc_hd__a211o_4
X_13370_ _13402_/A _19119_/A VGND VGND VPWR VPWR _13370_/X sky130_fd_sc_hd__or2_4
XANTENNA__12250__B1 _12249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25356_ _25356_/CLK _12977_/X HRESETn VGND VGND VPWR VPWR _25356_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22568_ _22549_/Y _22555_/Y _22564_/Y _21437_/X _22567_/X VGND VGND VPWR VPWR _22568_/X
+ sky130_fd_sc_hd__a32o_4
X_12321_ _24831_/Q VGND VGND VPWR VPWR _12321_/Y sky130_fd_sc_hd__inv_2
X_24307_ _24305_/CLK _24307_/D HRESETn VGND VGND VPWR VPWR _17515_/A sky130_fd_sc_hd__dfrtp_4
X_21519_ _24774_/Q _21519_/B VGND VGND VPWR VPWR _21519_/X sky130_fd_sc_hd__or2_4
XFILLER_103_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25287_ _25461_/CLK _25287_/D HRESETn VGND VGND VPWR VPWR _25287_/Q sky130_fd_sc_hd__dfrtp_4
X_22499_ _16246_/Y _22444_/A _15112_/Y _22441_/A VGND VGND VPWR VPWR _22500_/B sky130_fd_sc_hd__o22a_4
XFILLER_6_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15040_ _15034_/X _15035_/X _15037_/X _15039_/X VGND VGND VPWR VPWR _15055_/B sky130_fd_sc_hd__or4_4
XFILLER_108_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18269__B1 _23342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12252_ _12252_/A VGND VGND VPWR VPWR _12252_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25346__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24238_ _23516_/CLK _17926_/X HRESETn VGND VGND VPWR VPWR _13541_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_79_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12183_ _25426_/Q _12181_/Y _12291_/A _23178_/A VGND VGND VPWR VPWR _12183_/X sky130_fd_sc_hd__a2bb2o_4
X_24169_ _24171_/CLK _24169_/D HRESETn VGND VGND VPWR VPWR _18409_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_134_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16991_ _24377_/Q VGND VGND VPWR VPWR _17034_/B sky130_fd_sc_hd__inv_2
XFILLER_27_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13502__B1 _11833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15942_ HWDATA[28] VGND VGND VPWR VPWR _15942_/X sky130_fd_sc_hd__buf_2
X_18730_ _18603_/X _18729_/Y VGND VGND VPWR VPWR _18730_/X sky130_fd_sc_hd__or2_4
XFILLER_114_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21576__B1 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18661_ _16616_/Y _18681_/A _16620_/A _18639_/Y VGND VGND VPWR VPWR _18661_/X sky130_fd_sc_hd__a2bb2o_4
X_15873_ _12759_/Y _15869_/X _11757_/X _15872_/X VGND VGND VPWR VPWR _15873_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24981__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18178__A _17928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14824_ _14824_/A VGND VGND VPWR VPWR _14824_/X sky130_fd_sc_hd__buf_2
X_17612_ _17612_/A _17618_/A VGND VGND VPWR VPWR _17616_/B sky130_fd_sc_hd__or2_4
XFILLER_76_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18592_ _18592_/A VGND VGND VPWR VPWR _18592_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24299__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24910__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17543_ _17543_/A VGND VGND VPWR VPWR _17543_/Y sky130_fd_sc_hd__inv_2
X_14755_ _14679_/A VGND VGND VPWR VPWR _21372_/A sky130_fd_sc_hd__inv_2
XANTENNA__24228__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11967_ _11647_/X _11967_/B _11967_/C _11967_/D VGND VGND VPWR VPWR _11967_/X sky130_fd_sc_hd__and4_4
XFILLER_45_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13706_ _13702_/B _13680_/X _13705_/X _13703_/X _13693_/A VGND VGND VPWR VPWR _13706_/X
+ sky130_fd_sc_hd__a32o_4
X_17474_ _17474_/A _17451_/Y _17461_/X _17473_/X VGND VGND VPWR VPWR _17474_/X sky130_fd_sc_hd__or4_4
XFILLER_44_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15558__A1 _15548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14686_ _14697_/A _14697_/B VGND VGND VPWR VPWR _14686_/Y sky130_fd_sc_hd__nor2_4
X_11898_ _11869_/B _11897_/Y _11893_/A VGND VGND VPWR VPWR _11898_/X sky130_fd_sc_hd__o21a_4
X_16425_ _24578_/Q VGND VGND VPWR VPWR _16425_/Y sky130_fd_sc_hd__inv_2
X_19213_ _19210_/Y _19211_/X _19212_/X _19211_/X VGND VGND VPWR VPWR _19213_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13637_ _13637_/A VGND VGND VPWR VPWR _13638_/A sky130_fd_sc_hd__inv_2
XFILLER_60_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12954__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19144_ _19130_/A VGND VGND VPWR VPWR _19144_/X sky130_fd_sc_hd__buf_2
X_16356_ _16280_/X VGND VGND VPWR VPWR _16356_/X sky130_fd_sc_hd__buf_2
XANTENNA__21051__B _21026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24065__D _20461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13568_ _13570_/A VGND VGND VPWR VPWR _13568_/X sky130_fd_sc_hd__buf_2
XANTENNA__16507__B1 _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18638__A1_N _24519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15307_ _15135_/Y _15336_/C _15307_/C _15306_/X VGND VGND VPWR VPWR _15325_/B sky130_fd_sc_hd__or4_4
XFILLER_34_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12519_ _12511_/X _12513_/X _12516_/X _12518_/X VGND VGND VPWR VPWR _12558_/A sky130_fd_sc_hd__or4_4
X_19075_ _13369_/B VGND VGND VPWR VPWR _19075_/Y sky130_fd_sc_hd__inv_2
X_16287_ _23247_/A VGND VGND VPWR VPWR _16287_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13499_ _12023_/Y _13498_/X _11825_/X _13498_/X VGND VGND VPWR VPWR _13499_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18026_ _18133_/A _18026_/B VGND VGND VPWR VPWR _18026_/X sky130_fd_sc_hd__or2_4
X_15238_ _15209_/C _15165_/B VGND VGND VPWR VPWR _15239_/B sky130_fd_sc_hd__or2_4
XANTENNA__23259__A _23085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17257__A _17257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25016__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15169_ _14888_/Y _15169_/B VGND VGND VPWR VPWR _15170_/C sky130_fd_sc_hd__or2_4
XFILLER_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19977_ _19977_/A VGND VGND VPWR VPWR _22238_/B sky130_fd_sc_hd__inv_2
XFILLER_45_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18928_ _18927_/Y _18925_/X _17421_/X _18925_/X VGND VGND VPWR VPWR _23907_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18432__B1 _16234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18859_ _18855_/X _18859_/B _18857_/X _18858_/X VGND VGND VPWR VPWR _18865_/C sky130_fd_sc_hd__or4_4
XFILLER_83_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_114_0_HCLK clkbuf_7_57_0_HCLK/X VGND VGND VPWR VPWR _24162_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__23308__A1 _21512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23308__B2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_177_0_HCLK clkbuf_7_88_0_HCLK/X VGND VGND VPWR VPWR _24278_/CLK sky130_fd_sc_hd__clkbuf_1
X_21870_ _22425_/A _21868_/X _22963_/A _21869_/X VGND VGND VPWR VPWR _21870_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21319__B1 _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24651__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20821_ _24030_/Q _21209_/A _13653_/B VGND VGND VPWR VPWR _20821_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23540_ _23394_/CLK _23540_/D VGND VGND VPWR VPWR _19970_/A sky130_fd_sc_hd__dfxtp_4
X_20752_ _20743_/X _20751_/X _15597_/A _20747_/X VGND VGND VPWR VPWR _24013_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16746__B1 _15729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20683_ _13122_/A _23997_/Q _13123_/B VGND VGND VPWR VPWR _20683_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23471_ _23581_/CLK _23471_/D VGND VGND VPWR VPWR _20160_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_17_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12864__A _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25210_ _25093_/CLK _25210_/D HRESETn VGND VGND VPWR VPWR _25210_/Q sky130_fd_sc_hd__dfrtp_4
X_22422_ _22421_/X VGND VGND VPWR VPWR _22422_/X sky130_fd_sc_hd__buf_2
XANTENNA__22295__A1 _24541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25141_ _25141_/CLK _14372_/X HRESETn VGND VGND VPWR VPWR _25141_/Q sky130_fd_sc_hd__dfrtp_4
X_22353_ _22050_/X _22353_/B VGND VGND VPWR VPWR _22353_/X sky130_fd_sc_hd__or2_4
X_21304_ _21277_/Y VGND VGND VPWR VPWR _21304_/X sky130_fd_sc_hd__buf_2
X_22284_ _24778_/Q _21073_/B VGND VGND VPWR VPWR _22284_/X sky130_fd_sc_hd__or2_4
X_25072_ _25070_/CLK _25072_/D HRESETn VGND VGND VPWR VPWR _13566_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20058__B1 _19794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21235_ _14680_/X _21235_/B VGND VGND VPWR VPWR _21235_/X sky130_fd_sc_hd__or2_4
XFILLER_102_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24023_ _24055_/CLK _24023_/D HRESETn VGND VGND VPWR VPWR _20790_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_117_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16071__A _24705_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16277__A2 _15993_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21166_ _24200_/Q VGND VGND VPWR VPWR _21186_/A sky130_fd_sc_hd__inv_2
XFILLER_85_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20073__A3 _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22801__A _23021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20117_ _20117_/A VGND VGND VPWR VPWR _20117_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_10_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21097_ _22419_/A VGND VGND VPWR VPWR _21098_/A sky130_fd_sc_hd__inv_2
XFILLER_24_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24739__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_73_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_73_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20048_ _20047_/Y _20045_/X _19780_/X _20045_/X VGND VGND VPWR VPWR _20048_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24925_ _24926_/CLK _15514_/X HRESETn VGND VGND VPWR VPWR _11728_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12870_ _12869_/X VGND VGND VPWR VPWR _12871_/B sky130_fd_sc_hd__inv_2
XFILLER_85_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24392__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24856_ _24865_/CLK _15746_/X HRESETn VGND VGND VPWR VPWR _24856_/Q sky130_fd_sc_hd__dfrtp_4
X_11821_ HWDATA[10] VGND VGND VPWR VPWR _11821_/X sky130_fd_sc_hd__buf_2
X_23807_ _23805_/CLK _19213_/X VGND VGND VPWR VPWR _19210_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24321__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24787_ _24832_/CLK _24787_/D HRESETn VGND VGND VPWR VPWR _24787_/Q sky130_fd_sc_hd__dfrtp_4
X_21999_ _21998_/X VGND VGND VPWR VPWR _21999_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ scl_oen_o_S4 _14534_/X _14535_/Y _14539_/Y VGND VGND VPWR VPWR _14540_/X
+ sky130_fd_sc_hd__o22a_4
XANTENNA__17630__A _17630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11748_/Y _11742_/X _11749_/X _11751_/X VGND VGND VPWR VPWR _25536_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23738_ _23718_/CLK _23738_/D VGND VGND VPWR VPWR _18033_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16737__B1 _16384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21152__A _15670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14468_/Y _14466_/X _14470_/X _14466_/X VGND VGND VPWR VPWR _25110_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _24214_/Q VGND VGND VPWR VPWR _11683_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12774__A _25362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23669_ _23689_/CLK _23669_/D VGND VGND VPWR VPWR _23669_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_70_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16209_/Y _16205_/X _15952_/X _16205_/X VGND VGND VPWR VPWR _16210_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _13454_/A _13422_/B _13421_/X VGND VGND VPWR VPWR _13422_/X sky130_fd_sc_hd__or3_4
XFILLER_122_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22286__A1 _21413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25408_ _25020_/CLK _25408_/D HRESETn VGND VGND VPWR VPWR _25408_/Q sky130_fd_sc_hd__dfrtp_4
X_17190_ _22402_/A _24335_/Q _16347_/Y _17349_/A VGND VGND VPWR VPWR _17191_/D sky130_fd_sc_hd__o22a_4
XANTENNA__25527__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16141_ _16140_/Y _16138_/X _15897_/X _16138_/X VGND VGND VPWR VPWR _24678_/D sky130_fd_sc_hd__a2bb2o_4
X_13353_ _13317_/A _23640_/Q VGND VGND VPWR VPWR _13354_/C sky130_fd_sc_hd__or2_4
XFILLER_122_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25339_ _24852_/CLK _13062_/X HRESETn VGND VGND VPWR VPWR _25339_/Q sky130_fd_sc_hd__dfrtp_4
X_12304_ _13057_/A _24823_/Q _12303_/A _24823_/Q VGND VGND VPWR VPWR _12313_/A sky130_fd_sc_hd__a2bb2o_4
X_16072_ _16071_/Y _16067_/X _15986_/X _16067_/X VGND VGND VPWR VPWR _16072_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15712__A1 _15548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13284_ _13421_/A _13282_/X _13283_/X VGND VGND VPWR VPWR _13284_/X sky130_fd_sc_hd__and3_4
X_15023_ _15023_/A VGND VGND VPWR VPWR _15023_/Y sky130_fd_sc_hd__inv_2
X_19900_ _21803_/B _19895_/X _19625_/X _19895_/X VGND VGND VPWR VPWR _23568_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12235_ _12235_/A VGND VGND VPWR VPWR _12235_/X sky130_fd_sc_hd__buf_2
XFILLER_108_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19831_ _23593_/Q VGND VGND VPWR VPWR _19831_/Y sky130_fd_sc_hd__inv_2
X_12166_ _12166_/A _18370_/B VGND VGND VPWR VPWR _12166_/X sky130_fd_sc_hd__and2_4
XFILLER_111_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18662__B1 _16547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19762_ _19761_/Y _19759_/X _19715_/X _19759_/X VGND VGND VPWR VPWR _19762_/X sky130_fd_sc_hd__a2bb2o_4
X_12097_ _12096_/X VGND VGND VPWR VPWR _12097_/X sky130_fd_sc_hd__buf_2
X_16974_ _24368_/Q VGND VGND VPWR VPWR _17038_/B sky130_fd_sc_hd__inv_2
X_18713_ _18705_/A _18711_/A VGND VGND VPWR VPWR _18713_/X sky130_fd_sc_hd__or2_4
XANTENNA__17217__B2 _17350_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15925_ _15777_/B _15925_/B VGND VGND VPWR VPWR _15925_/X sky130_fd_sc_hd__or2_4
X_19693_ _19692_/Y _19690_/X _19547_/X _19690_/X VGND VGND VPWR VPWR _19693_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24409__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11853__A _16359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15856_ _15894_/A VGND VGND VPWR VPWR _15857_/A sky130_fd_sc_hd__buf_2
X_18644_ _16587_/Y _18688_/A _16587_/Y _18688_/A VGND VGND VPWR VPWR _18645_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14807_ _14807_/A _14807_/B _14807_/C VGND VGND VPWR VPWR _14807_/X sky130_fd_sc_hd__or3_4
XFILLER_18_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24062__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15787_ _15819_/A VGND VGND VPWR VPWR _15795_/A sky130_fd_sc_hd__buf_2
X_18575_ _18411_/Y _18575_/B VGND VGND VPWR VPWR _18575_/Y sky130_fd_sc_hd__nand2_4
X_12999_ _13029_/A _12999_/B _12999_/C _12999_/D VGND VGND VPWR VPWR _12999_/X sky130_fd_sc_hd__or4_4
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14738_ _14726_/X _14730_/Y VGND VGND VPWR VPWR _14738_/Y sky130_fd_sc_hd__nor2_4
X_17526_ _25524_/Q _17525_/Y _11840_/Y _24283_/Q VGND VGND VPWR VPWR _17526_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21062__A _15784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17457_ _17457_/A VGND VGND VPWR VPWR _17457_/Y sky130_fd_sc_hd__inv_2
X_14669_ _25059_/Q VGND VGND VPWR VPWR _19152_/A sky130_fd_sc_hd__buf_2
X_16408_ HWDATA[18] VGND VGND VPWR VPWR _16408_/X sky130_fd_sc_hd__buf_2
XFILLER_32_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25268__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17388_ _23969_/Q _17388_/B VGND VGND VPWR VPWR _17388_/X sky130_fd_sc_hd__or2_4
XFILLER_20_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16339_ _24609_/Q VGND VGND VPWR VPWR _16339_/Y sky130_fd_sc_hd__inv_2
X_19127_ _25059_/Q _13613_/X _14659_/A VGND VGND VPWR VPWR _19399_/C sky130_fd_sc_hd__or3_4
XFILLER_12_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19058_ _23861_/Q VGND VGND VPWR VPWR _19058_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18009_ _18150_/A _19132_/A VGND VGND VPWR VPWR _18012_/B sky130_fd_sc_hd__or2_4
XANTENNA__18248__A3 _18247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21020_ _22929_/A VGND VGND VPWR VPWR _22523_/A sky130_fd_sc_hd__buf_2
XFILLER_86_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18653__B1 _16597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17715__A _21192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24832__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22971_ _22971_/A _22898_/X VGND VGND VPWR VPWR _22971_/X sky130_fd_sc_hd__or2_4
XANTENNA__12859__A _12859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14690__B2 _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24710_ _24712_/CLK _16058_/X HRESETn VGND VGND VPWR VPWR _24710_/Q sky130_fd_sc_hd__dfrtp_4
X_21922_ _21916_/X _21921_/X _17722_/A VGND VGND VPWR VPWR _21922_/X sky130_fd_sc_hd__o21a_4
XFILLER_67_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20763__A1 _13119_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24641_ _24162_/CLK _16252_/X HRESETn VGND VGND VPWR VPWR _22294_/A sky130_fd_sc_hd__dfrtp_4
X_21853_ _24707_/Q _22406_/B _21103_/A _21852_/X VGND VGND VPWR VPWR _21854_/C sky130_fd_sc_hd__a211o_4
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20804_ _20804_/A _20799_/A _13136_/X VGND VGND VPWR VPWR _20804_/X sky130_fd_sc_hd__or3_4
XANTENNA__17450__A _17449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24572_ _24572_/CLK _16435_/X HRESETn VGND VGND VPWR VPWR _15126_/A sky130_fd_sc_hd__dfrtp_4
X_21784_ _21777_/Y _21783_/Y _13784_/C VGND VGND VPWR VPWR _21784_/X sky130_fd_sc_hd__o21a_4
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23523_ _23394_/CLK _23523_/D VGND VGND VPWR VPWR _20026_/A sky130_fd_sc_hd__dfxtp_4
X_20735_ _13133_/A _13133_/B VGND VGND VPWR VPWR _20740_/B sky130_fd_sc_hd__or2_4
XFILLER_24_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16066__A _24707_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23454_ _23478_/CLK _23454_/D VGND VGND VPWR VPWR _20205_/A sky130_fd_sc_hd__dfxtp_4
X_20666_ _14281_/X VGND VGND VPWR VPWR _20666_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21122__D _13813_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22405_ _22658_/A _22405_/B VGND VGND VPWR VPWR _22417_/C sky130_fd_sc_hd__nor2_4
XANTENNA__21700__A _21108_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20597_ _25096_/Q _20594_/Y _20595_/Y _14495_/X _20596_/X VGND VGND VPWR VPWR _20597_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_52_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23385_ _23384_/CLK _23385_/D VGND VGND VPWR VPWR _23385_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18281__A _17702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22515__B _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25124_ _24364_/CLK _25124_/D HRESETn VGND VGND VPWR VPWR _25124_/Q sky130_fd_sc_hd__dfstp_4
X_22336_ _21945_/A _19929_/Y VGND VGND VPWR VPWR _22337_/C sky130_fd_sc_hd__or2_4
XANTENNA__23217__B1 _24731_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25055_ _25055_/CLK _14737_/X HRESETn VGND VGND VPWR VPWR _25055_/Q sky130_fd_sc_hd__dfrtp_4
X_22267_ _22267_/A _22266_/X VGND VGND VPWR VPWR _22267_/X sky130_fd_sc_hd__or2_4
XANTENNA__18239__A3 _11803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12020_ _12020_/A VGND VGND VPWR VPWR _12020_/Y sky130_fd_sc_hd__inv_2
X_24006_ _24035_/CLK _20720_/Y HRESETn VGND VGND VPWR VPWR _20717_/A sky130_fd_sc_hd__dfrtp_4
X_21218_ _25286_/Q _21112_/B VGND VGND VPWR VPWR _21218_/Y sky130_fd_sc_hd__nor2_4
XFILLER_133_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18644__B1 _16587_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22198_ _21240_/X _19913_/Y VGND VGND VPWR VPWR _22198_/X sky130_fd_sc_hd__or2_4
XFILLER_133_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17625__A _17557_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21149_ _16622_/Y _21154_/B VGND VGND VPWR VPWR _21149_/X sky130_fd_sc_hd__or2_4
XANTENNA__24573__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14690__A2_N _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14130__B1 _14128_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13971_ _13971_/A VGND VGND VPWR VPWR _13971_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24502__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23065__C _23064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15710_ _15740_/A VGND VGND VPWR VPWR _15711_/A sky130_fd_sc_hd__buf_2
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12922_ _12753_/X _12903_/X _12874_/X _12919_/Y VGND VGND VPWR VPWR _12922_/X sky130_fd_sc_hd__a211o_4
XFILLER_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24908_ _24025_/CLK _24908_/D HRESETn VGND VGND VPWR VPWR _24908_/Q sky130_fd_sc_hd__dfrtp_4
X_16690_ _24478_/Q VGND VGND VPWR VPWR _22634_/A sky130_fd_sc_hd__inv_2
XFILLER_59_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21951__B1 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16995__A1_N _24704_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15641_ _15641_/A VGND VGND VPWR VPWR _22824_/A sky130_fd_sc_hd__buf_2
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23362__A _21005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12853_ _12887_/A _12886_/A _12841_/X _12852_/X VGND VGND VPWR VPWR _12854_/B sky130_fd_sc_hd__or4_4
Xclkbuf_8_160_0_HCLK clkbuf_7_80_0_HCLK/X VGND VGND VPWR VPWR _25497_/CLK sky130_fd_sc_hd__clkbuf_1
X_24839_ _24840_/CLK _15780_/X HRESETn VGND VGND VPWR VPWR _24839_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_3_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_92_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15630__B1 _15471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11804_ _11803_/X VGND VGND VPWR VPWR _11804_/X sky130_fd_sc_hd__buf_2
X_18360_ _18359_/Y _17478_/X _18359_/A _17482_/X VGND VGND VPWR VPWR _18361_/A sky130_fd_sc_hd__o22a_4
XFILLER_15_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15572_ _15572_/A VGND VGND VPWR VPWR _15572_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_17_0_HCLK clkbuf_7_8_0_HCLK/X VGND VGND VPWR VPWR _25141_/CLK sky130_fd_sc_hd__clkbuf_1
X_12784_ _12954_/A VGND VGND VPWR VPWR _12955_/A sky130_fd_sc_hd__inv_2
XFILLER_61_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21703__B1 _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17311_ _17311_/A VGND VGND VPWR VPWR _17311_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14521_/X _14522_/X _14480_/A _14517_/X VGND VGND VPWR VPWR _14523_/X sky130_fd_sc_hd__o22a_4
XPHY_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11735_ _21314_/A VGND VGND VPWR VPWR _21018_/A sky130_fd_sc_hd__buf_2
X_18291_ _24201_/Q VGND VGND VPWR VPWR _18291_/X sky130_fd_sc_hd__buf_2
XPHY_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17242_/A VGND VGND VPWR VPWR _17243_/D sky130_fd_sc_hd__inv_2
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _14453_/Y VGND VGND VPWR VPWR _14454_/X sky130_fd_sc_hd__buf_2
XANTENNA__25361__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11658_/X _11666_/B _11662_/X _11666_/D VGND VGND VPWR VPWR _11666_/X sky130_fd_sc_hd__or4_4
XFILLER_70_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22706__A _22706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _13270_/A _23438_/Q VGND VGND VPWR VPWR _13405_/X sky130_fd_sc_hd__or2_4
XANTENNA__21610__A _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17173_ _16322_/Y _24344_/Q _16322_/Y _24344_/Q VGND VGND VPWR VPWR _17173_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14385_ _20496_/C _14382_/X _13835_/X _14384_/X VGND VGND VPWR VPWR _14385_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16124_ _22774_/A VGND VGND VPWR VPWR _16124_/Y sky130_fd_sc_hd__inv_2
X_13336_ _24190_/Q VGND VGND VPWR VPWR _17452_/B sky130_fd_sc_hd__buf_2
XFILLER_116_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16055_ _16054_/Y _16052_/X _15758_/X _16052_/X VGND VGND VPWR VPWR _16055_/X sky130_fd_sc_hd__a2bb2o_4
X_13267_ _13457_/A _13265_/X _13267_/C VGND VGND VPWR VPWR _13267_/X sky130_fd_sc_hd__and3_4
XFILLER_29_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15006_ _15179_/A _15005_/A _15180_/A _15005_/Y VGND VGND VPWR VPWR _15012_/B sky130_fd_sc_hd__o22a_4
XFILLER_68_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12218_ _12399_/A _24764_/Q _12385_/A _12217_/Y VGND VGND VPWR VPWR _12218_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22431__A1 _12769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13198_ _13196_/Y VGND VGND VPWR VPWR _13198_/X sky130_fd_sc_hd__buf_2
XFILLER_69_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22431__B2 _21413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19814_ _23599_/Q VGND VGND VPWR VPWR _19814_/Y sky130_fd_sc_hd__inv_2
X_12149_ _24100_/Q _12147_/B _12148_/Y VGND VGND VPWR VPWR _12149_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23256__B _23082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19745_ _23622_/Q VGND VGND VPWR VPWR _19745_/Y sky130_fd_sc_hd__inv_2
X_16957_ _21004_/B _16955_/X _16956_/Y VGND VGND VPWR VPWR _24392_/D sky130_fd_sc_hd__o21a_4
XANTENNA__24243__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22734__A2 _22525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15908_ _12788_/Y _15904_/X _15477_/X _15904_/X VGND VGND VPWR VPWR _24774_/D sky130_fd_sc_hd__a2bb2o_4
X_19676_ _19676_/A VGND VGND VPWR VPWR _19676_/X sky130_fd_sc_hd__buf_2
XANTENNA__16949__B1 _16156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16888_ _19797_/A VGND VGND VPWR VPWR _16888_/X sky130_fd_sc_hd__buf_2
X_18627_ _24521_/Q _24132_/Q _16574_/Y _18626_/Y VGND VGND VPWR VPWR _18635_/A sky130_fd_sc_hd__o22a_4
XFILLER_37_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15839_ _12334_/Y _15833_/X _15477_/X _15833_/X VGND VGND VPWR VPWR _24809_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15621__B1 _15620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25449__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18558_ _16448_/A _18475_/D VGND VGND VPWR VPWR _18592_/A sky130_fd_sc_hd__or2_4
XANTENNA__21504__B _21504_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17701__C _21686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17509_ _11828_/A _24286_/Q _11828_/Y _17676_/A VGND VGND VPWR VPWR _17509_/X sky130_fd_sc_hd__o22a_4
X_18489_ _18489_/A VGND VGND VPWR VPWR _18489_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17374__B1 _17289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12845__C _12976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20520_ _24068_/Q _20519_/X _20508_/X VGND VGND VPWR VPWR _20520_/X sky130_fd_sc_hd__a21o_4
XFILLER_53_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15385__C1 _15339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20451_ _20451_/A _20449_/Y VGND VGND VPWR VPWR _24080_/D sky130_fd_sc_hd__or2_4
XFILLER_20_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21520__A _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25031__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20382_ _20317_/X _20379_/X _13835_/A _22390_/A _20381_/X VGND VGND VPWR VPWR _23387_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22670__A1 _16234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23170_ _23170_/A VGND VGND VPWR VPWR _23207_/A sky130_fd_sc_hd__buf_2
X_22121_ _24777_/Q _21530_/X VGND VGND VPWR VPWR _22121_/X sky130_fd_sc_hd__or2_4
XFILLER_12_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22052_ _21887_/X _19248_/Y VGND VGND VPWR VPWR _22052_/X sky130_fd_sc_hd__or2_4
XFILLER_133_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21003_ _21003_/A _21091_/A VGND VGND VPWR VPWR _21003_/X sky130_fd_sc_hd__and2_4
XANTENNA__13973__A _20490_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12910__A1 _12849_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25122__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22954_ _12257_/Y _22268_/X _22712_/X _12366_/Y _22840_/X VGND VGND VPWR VPWR _22955_/B
+ sky130_fd_sc_hd__o32a_4
XANTENNA__25185__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21905_ _21601_/A _21903_/X _21905_/C VGND VGND VPWR VPWR _21905_/X sky130_fd_sc_hd__and3_4
XFILLER_55_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22885_ _22885_/A VGND VGND VPWR VPWR _22885_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_233_0_HCLK clkbuf_8_233_0_HCLK/A VGND VGND VPWR VPWR _24780_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__23588__CLK _23498_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24624_ _24356_/CLK _24624_/D HRESETn VGND VGND VPWR VPWR _24624_/Q sky130_fd_sc_hd__dfrtp_4
X_21836_ _21836_/A _22927_/A VGND VGND VPWR VPWR _21836_/X sky130_fd_sc_hd__or2_4
XANTENNA__12426__B1 _12252_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21414__B _21073_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24555_ _24555_/CLK _16487_/X HRESETn VGND VGND VPWR VPWR _16485_/A sky130_fd_sc_hd__dfrtp_4
X_21767_ _21233_/X VGND VGND VPWR VPWR _21767_/X sky130_fd_sc_hd__buf_2
XFILLER_52_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13213__A _13227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23506_ _24208_/CLK _23506_/D VGND VGND VPWR VPWR _13273_/B sky130_fd_sc_hd__dfxtp_4
X_20718_ _20717_/Y _20713_/X _13130_/B VGND VGND VPWR VPWR _20718_/X sky130_fd_sc_hd__o21a_4
XFILLER_12_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24486_ _24447_/CLK _24486_/D HRESETn VGND VGND VPWR VPWR _24486_/Q sky130_fd_sc_hd__dfrtp_4
X_21698_ _16640_/A _21697_/X _21427_/X _24810_/Q _21323_/X VGND VGND VPWR VPWR _21699_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22526__A _22798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23437_ _23904_/CLK _23437_/D VGND VGND VPWR VPWR _23437_/Q sky130_fd_sc_hd__dfxtp_4
X_20649_ _20648_/X VGND VGND VPWR VPWR _23978_/D sky130_fd_sc_hd__inv_2
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22110__B1 _22109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14170_ _14098_/A VGND VGND VPWR VPWR _14170_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22661__A1 _12430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23368_ _24026_/CLK _20674_/A VGND VGND VPWR VPWR _13140_/A sky130_fd_sc_hd__dfxtp_4
X_13121_ _23999_/Q VGND VGND VPWR VPWR _13121_/Y sky130_fd_sc_hd__inv_2
X_25107_ _24945_/CLK _14479_/X HRESETn VGND VGND VPWR VPWR _25107_/Q sky130_fd_sc_hd__dfrtp_4
X_22319_ _14807_/A _21549_/B _20663_/A _22172_/B VGND VGND VPWR VPWR _22319_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24754__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23299_ _23208_/A _23299_/B _23299_/C _23299_/D VGND VGND VPWR VPWR _23299_/X sky130_fd_sc_hd__or4_4
X_13052_ _12349_/Y _13052_/B VGND VGND VPWR VPWR _13052_/X sky130_fd_sc_hd__or2_4
XANTENNA__23357__A _23344_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25038_ _25029_/CLK _25038_/D HRESETn VGND VGND VPWR VPWR _14802_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24324__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12003_ _13509_/A _11991_/A _13509_/A _11991_/A VGND VGND VPWR VPWR _12003_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17355__A _17350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17860_ _17862_/B VGND VGND VPWR VPWR _17861_/B sky130_fd_sc_hd__inv_2
X_16811_ _16807_/A VGND VGND VPWR VPWR _16811_/X sky130_fd_sc_hd__buf_2
XFILLER_78_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17791_ _17791_/A VGND VGND VPWR VPWR _17791_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12499__A _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22177__B1 _23962_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19530_ _23694_/Q VGND VGND VPWR VPWR _19530_/Y sky130_fd_sc_hd__inv_2
X_13954_ _13899_/X _13901_/X _13905_/C _13904_/Y VGND VGND VPWR VPWR _13954_/X sky130_fd_sc_hd__or4_4
X_16742_ _16741_/Y _16739_/X _15725_/X _16739_/X VGND VGND VPWR VPWR _16742_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_43_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_87_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12905_ _12849_/D _12905_/B VGND VGND VPWR VPWR _12905_/X sky130_fd_sc_hd__or2_4
X_16673_ _24485_/Q VGND VGND VPWR VPWR _16673_/Y sky130_fd_sc_hd__inv_2
X_19461_ _19461_/A VGND VGND VPWR VPWR _19461_/Y sky130_fd_sc_hd__inv_2
X_13885_ _20467_/A VGND VGND VPWR VPWR _20490_/A sky130_fd_sc_hd__buf_2
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15603__B1 _11804_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18412_ _22294_/A _24152_/Q _16251_/Y _18411_/Y VGND VGND VPWR VPWR _18412_/X sky130_fd_sc_hd__o22a_4
X_12836_ _12836_/A _12815_/X _12827_/X _12836_/D VGND VGND VPWR VPWR _12836_/X sky130_fd_sc_hd__or4_4
X_15624_ _22281_/A _15617_/X _15623_/X _15617_/X VGND VGND VPWR VPWR _24886_/D sky130_fd_sc_hd__a2bb2o_4
X_19392_ _19384_/A VGND VGND VPWR VPWR _19392_/X sky130_fd_sc_hd__buf_2
XFILLER_62_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12968__A1 _12819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15555_ _21154_/B VGND VGND VPWR VPWR _22695_/B sky130_fd_sc_hd__buf_2
X_18343_ _13174_/X _18345_/A _18340_/X VGND VGND VPWR VPWR _24192_/D sky130_fd_sc_hd__o21a_4
XANTENNA__22139__C _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12767_ _25363_/Q VGND VGND VPWR VPWR _12846_/B sky130_fd_sc_hd__inv_2
XANTENNA__14219__A _14219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17356__B1 _17289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _23951_/Q VGND VGND VPWR VPWR _14517_/A sky130_fd_sc_hd__inv_2
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _15549_/A _12052_/B VGND VGND VPWR VPWR _15991_/D sky130_fd_sc_hd__or2_4
X_18274_ _17729_/A VGND VGND VPWR VPWR _18275_/A sky130_fd_sc_hd__buf_2
X_15486_ _15484_/A _15484_/B _15485_/Y _14553_/Y VGND VGND VPWR VPWR _15486_/X sky130_fd_sc_hd__a211o_4
X_12698_ _12698_/A _12696_/X _12697_/X VGND VGND VPWR VPWR _25401_/D sky130_fd_sc_hd__and3_4
XANTENNA__15906__B2 _15864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14437_ _14436_/Y VGND VGND VPWR VPWR _14437_/X sky130_fd_sc_hd__buf_2
X_17225_ _16358_/Y _24331_/Q _24600_/Q _17206_/X VGND VGND VPWR VPWR _17229_/A sky130_fd_sc_hd__a2bb2o_4
X_11649_ _17481_/C VGND VGND VPWR VPWR _21504_/A sky130_fd_sc_hd__buf_2
XFILLER_122_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17156_ _17156_/A _17160_/A VGND VGND VPWR VPWR _17156_/Y sky130_fd_sc_hd__nand2_4
X_14368_ _25143_/Q _14348_/Y _25142_/Q _14344_/X VGND VGND VPWR VPWR _14368_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22652__A1 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18856__B1 _24558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22652__B2 _21533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16107_ _16105_/Y _16101_/X _15949_/X _16106_/X VGND VGND VPWR VPWR _24692_/D sky130_fd_sc_hd__a2bb2o_4
X_13319_ _13387_/A _13319_/B VGND VGND VPWR VPWR _13319_/X sky130_fd_sc_hd__or2_4
X_17087_ _17048_/D _17065_/X _17048_/B VGND VGND VPWR VPWR _17087_/X sky130_fd_sc_hd__o21a_4
X_14299_ _14299_/A VGND VGND VPWR VPWR _14299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24495__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16038_ _16037_/Y _16035_/X _11800_/X _16035_/X VGND VGND VPWR VPWR _16038_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24424__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20415__B1 _18267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_125_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_125_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17265__A _17264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16095__B1 _15940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17989_ _18211_/A _17989_/B VGND VGND VPWR VPWR _17992_/B sky130_fd_sc_hd__or2_4
XFILLER_42_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15842__B1 _24807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24109__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19728_ _19728_/A _17462_/Y _18333_/X _18335_/X VGND VGND VPWR VPWR _19729_/A sky130_fd_sc_hd__or4_4
XANTENNA__19033__B1 _18940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12202__A _12202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19659_ _19657_/Y _19653_/X _19658_/X _19638_/Y VGND VGND VPWR VPWR _19659_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25283__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22670_ _16234_/Y _22444_/X _16421_/Y _22441_/X VGND VGND VPWR VPWR _22671_/B sky130_fd_sc_hd__o22a_4
XFILLER_0_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21621_ _21616_/A _19858_/Y VGND VGND VPWR VPWR _21621_/X sky130_fd_sc_hd__or2_4
XANTENNA__25212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_63_0_HCLK clkbuf_8_63_0_HCLK/A VGND VGND VPWR VPWR _24345_/CLK sky130_fd_sc_hd__clkbuf_1
X_24340_ _24612_/CLK _17343_/Y HRESETn VGND VGND VPWR VPWR _24340_/Q sky130_fd_sc_hd__dfrtp_4
X_21552_ _21552_/A VGND VGND VPWR VPWR _21552_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22346__A _21455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20503_ _24070_/Q _20503_/B VGND VGND VPWR VPWR _20504_/C sky130_fd_sc_hd__and2_4
XFILLER_138_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24271_ _24267_/CLK _17791_/Y HRESETn VGND VGND VPWR VPWR _17740_/A sky130_fd_sc_hd__dfrtp_4
X_21483_ _21449_/A _21483_/B VGND VGND VPWR VPWR _21485_/B sky130_fd_sc_hd__or2_4
XANTENNA__12872__A _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23222_ _23281_/A _23222_/B _23222_/C _23221_/X VGND VGND VPWR VPWR _23222_/X sky130_fd_sc_hd__or4_4
X_20434_ _20443_/A _20433_/X VGND VGND VPWR VPWR _20458_/A sky130_fd_sc_hd__and2_4
XANTENNA__13687__B _13686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18847__B1 _24540_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23153_ _22975_/X _23152_/X _23044_/X _25533_/Q _23111_/X VGND VGND VPWR VPWR _23153_/X
+ sky130_fd_sc_hd__a32o_4
X_20365_ _23393_/Q VGND VGND VPWR VPWR _22027_/B sky130_fd_sc_hd__inv_2
X_22104_ _12959_/A _21009_/X _20837_/Y _22103_/X VGND VGND VPWR VPWR _22104_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15676__A3 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20296_ _23419_/Q VGND VGND VPWR VPWR _22347_/B sky130_fd_sc_hd__inv_2
XANTENNA__24165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23084_ _14919_/A _22833_/X _22090_/X _23083_/X VGND VGND VPWR VPWR _23085_/C sky130_fd_sc_hd__a211o_4
XANTENNA__20406__B1 _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22946__A2 _22790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22035_ _22035_/A _22034_/X VGND VGND VPWR VPWR _22035_/X sky130_fd_sc_hd__and2_4
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19024__B1 _18997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23986_ _23964_/CLK _23985_/Q HRESETn VGND VGND VPWR VPWR _23986_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21425__A _21525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22937_ _24522_/Q _22393_/X _15668_/A _22936_/X VGND VGND VPWR VPWR _22938_/C sky130_fd_sc_hd__a211o_4
XFILLER_21_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13670_ _13670_/A _13669_/Y VGND VGND VPWR VPWR _13670_/X sky130_fd_sc_hd__and2_4
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12370__A2_N _12368_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22868_ _22778_/A _22856_/X _22868_/C _22867_/X VGND VGND VPWR VPWR _22868_/X sky130_fd_sc_hd__or4_4
X_12621_ _12524_/Y _12620_/X VGND VGND VPWR VPWR _12642_/B sky130_fd_sc_hd__or2_4
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24607_ _24606_/CLK _16346_/X HRESETn VGND VGND VPWR VPWR _16345_/A sky130_fd_sc_hd__dfrtp_4
X_21819_ _21994_/A _21818_/X _24216_/Q _13815_/X VGND VGND VPWR VPWR _21819_/X sky130_fd_sc_hd__o22a_4
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21134__B2 _12059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22331__B1 _17722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22799_ _15003_/A _22654_/X _22798_/X VGND VGND VPWR VPWR _22799_/X sky130_fd_sc_hd__o21a_4
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15340_ _15080_/Y _15338_/X _15339_/X VGND VGND VPWR VPWR _15340_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_12_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12552_ _12552_/A VGND VGND VPWR VPWR _12552_/Y sky130_fd_sc_hd__inv_2
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24538_ _24545_/CLK _16532_/X HRESETn VGND VGND VPWR VPWR _21837_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22256__A _21681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21160__A _17447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15271_ _15282_/A _15267_/X _15271_/C VGND VGND VPWR VPWR _15271_/X sky130_fd_sc_hd__and3_4
XFILLER_36_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ _12220_/X _12481_/A VGND VGND VPWR VPWR _12483_/X sky130_fd_sc_hd__or2_4
XFILLER_89_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24469_ _24033_/CLK _16713_/X HRESETn VGND VGND VPWR VPWR _16711_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24935__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17010_ _24725_/Q _17048_/B _16024_/Y _17007_/A VGND VGND VPWR VPWR _17010_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222_ _14195_/A VGND VGND VPWR VPWR _14223_/B sky130_fd_sc_hd__buf_2
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13597__B _14433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14153_ _14115_/A _14115_/B _14115_/A _14115_/B VGND VGND VPWR VPWR _14154_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA_clkbuf_5_27_0_HCLK_A clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13104_ _12363_/Y _13081_/B _13101_/Y _13031_/X VGND VGND VPWR VPWR _13105_/A sky130_fd_sc_hd__a211o_4
XFILLER_113_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22703__B _21511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14084_ _14084_/A VGND VGND VPWR VPWR _14084_/X sky130_fd_sc_hd__buf_2
X_18961_ _16442_/A VGND VGND VPWR VPWR _18961_/X sky130_fd_sc_hd__buf_2
XANTENNA__20504__A _20490_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22398__B1 _23314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13035_ _13038_/A _13035_/B _13034_/Y VGND VGND VPWR VPWR _13035_/X sky130_fd_sc_hd__and3_4
X_17912_ _13590_/A _14769_/X _14620_/A VGND VGND VPWR VPWR _17912_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22937__A2 _22393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18892_ _18868_/Y _18882_/Y _23946_/Q _24106_/Q _20582_/B VGND VGND VPWR VPWR _24106_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_67_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17843_ _17753_/Y _17837_/X _17790_/A _17840_/B VGND VGND VPWR VPWR _17844_/A sky130_fd_sc_hd__a211o_4
XFILLER_39_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17540__A1_N _11844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17774_ _17774_/A VGND VGND VPWR VPWR _17774_/Y sky130_fd_sc_hd__inv_2
X_14986_ _14986_/A VGND VGND VPWR VPWR _15199_/A sky130_fd_sc_hd__inv_2
X_19513_ _19513_/A VGND VGND VPWR VPWR _22340_/B sky130_fd_sc_hd__inv_2
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16725_ _16725_/A _16725_/B _22574_/A _21314_/B VGND VGND VPWR VPWR _16725_/X sky130_fd_sc_hd__and4_4
XANTENNA__21335__A _21335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13937_ _13921_/Y VGND VGND VPWR VPWR _13952_/A sky130_fd_sc_hd__buf_2
XANTENNA__24082__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11861__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19444_ _23724_/Q VGND VGND VPWR VPWR _19444_/Y sky130_fd_sc_hd__inv_2
X_13868_ _13852_/X _13866_/X _14254_/A _13867_/X VGND VGND VPWR VPWR _13868_/X sky130_fd_sc_hd__o22a_4
X_16656_ _16655_/Y _16651_/X _16297_/X _16651_/X VGND VGND VPWR VPWR _16656_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12819_ _12819_/A VGND VGND VPWR VPWR _12819_/X sky130_fd_sc_hd__buf_2
X_15607_ _24892_/Q VGND VGND VPWR VPWR _15607_/Y sky130_fd_sc_hd__inv_2
X_19375_ _19374_/Y _19369_/X _19307_/X _19355_/Y VGND VGND VPWR VPWR _23749_/D sky130_fd_sc_hd__a2bb2o_4
X_13799_ _13799_/A VGND VGND VPWR VPWR _13799_/Y sky130_fd_sc_hd__inv_2
X_16587_ _16587_/A VGND VGND VPWR VPWR _16587_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20893__B _20884_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18326_ _18325_/X VGND VGND VPWR VPWR _18326_/X sky130_fd_sc_hd__buf_2
X_15538_ _15535_/A VGND VGND VPWR VPWR _15538_/X sky130_fd_sc_hd__buf_2
XANTENNA__21070__A _23019_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15469_ _15467_/Y _15463_/X _14418_/X _15468_/X VGND VGND VPWR VPWR _15469_/X sky130_fd_sc_hd__a2bb2o_4
X_18257_ _11683_/Y _18233_/A _16717_/X _18233_/A VGND VGND VPWR VPWR _18257_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24676__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17208_ _24600_/Q _17206_/X _16352_/A _17365_/A VGND VGND VPWR VPWR _17211_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18829__B1 _16476_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18188_ _18220_/A _18188_/B _18188_/C VGND VGND VPWR VPWR _18192_/B sky130_fd_sc_hd__and3_4
XFILLER_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24605__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17139_ _17143_/A _17135_/X _17138_/Y VGND VGND VPWR VPWR _24370_/D sky130_fd_sc_hd__and3_4
XANTENNA__22613__B _22613_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20150_ _20146_/Y _20149_/X _20079_/X _20149_/X VGND VGND VPWR VPWR _23476_/D sky130_fd_sc_hd__a2bb2o_4
X_20081_ _23499_/Q VGND VGND VPWR VPWR _22194_/B sky130_fd_sc_hd__inv_2
XANTENNA__16068__B1 _15471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15815__B1 _11791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19006__B1 _18961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23840_ _23854_/CLK _19118_/X VGND VGND VPWR VPWR _13338_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__25464__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19519__A2_N _19516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23771_ _23772_/CLK _23771_/D VGND VGND VPWR VPWR _17974_/B sky130_fd_sc_hd__dfxtp_4
X_20983_ sda_oen_o_S4 _25086_/Q _20978_/A _14037_/X _20982_/Y VGND VGND VPWR VPWR
+ _23923_/D sky130_fd_sc_hd__a32o_4
XANTENNA__11771__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25510_ _25508_/CLK _25510_/D HRESETn VGND VGND VPWR VPWR _25510_/Q sky130_fd_sc_hd__dfrtp_4
X_22722_ _24582_/Q _22722_/B VGND VGND VPWR VPWR _22722_/X sky130_fd_sc_hd__or2_4
XFILLER_129_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25441_ _25425_/CLK _25441_/D HRESETn VGND VGND VPWR VPWR _12284_/A sky130_fd_sc_hd__dfrtp_4
X_22653_ _22653_/A VGND VGND VPWR VPWR _22653_/Y sky130_fd_sc_hd__inv_2
X_21604_ _21630_/A _20202_/Y VGND VGND VPWR VPWR _21605_/C sky130_fd_sc_hd__or2_4
X_25372_ _25374_/CLK _25372_/D HRESETn VGND VGND VPWR VPWR _12810_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22584_ _16510_/A _22422_/X _22527_/X VGND VGND VPWR VPWR _22584_/X sky130_fd_sc_hd__o21a_4
XFILLER_107_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24323_ _23967_/CLK _24323_/D HRESETn VGND VGND VPWR VPWR _24323_/Q sky130_fd_sc_hd__dfstp_4
X_21535_ _21524_/X _21528_/Y _22705_/A _21534_/X VGND VGND VPWR VPWR _21535_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22616__A1 _17249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24254_ _24673_/CLK _17863_/X HRESETn VGND VGND VPWR VPWR _16918_/A sky130_fd_sc_hd__dfrtp_4
X_21466_ _21658_/A _19945_/Y VGND VGND VPWR VPWR _21467_/C sky130_fd_sc_hd__or2_4
XANTENNA__24346__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_7_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23205_ _15015_/A _22998_/X _23172_/X VGND VGND VPWR VPWR _23205_/X sky130_fd_sc_hd__o21a_4
X_20417_ _20416_/Y _20412_/X _15647_/X _20399_/Y VGND VGND VPWR VPWR _23371_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22092__A2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24185_ _24373_/CLK _24185_/D HRESETn VGND VGND VPWR VPWR _18369_/A sky130_fd_sc_hd__dfrtp_4
X_21397_ _21385_/A _20059_/Y VGND VGND VPWR VPWR _21397_/X sky130_fd_sc_hd__or2_4
XANTENNA__16802__A _16807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12107__A _12119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23136_ _16809_/A _22929_/X _22997_/X _23135_/X VGND VGND VPWR VPWR _23136_/X sky130_fd_sc_hd__a211o_4
X_20348_ _20347_/Y _20345_/X _19622_/A _20345_/X VGND VGND VPWR VPWR _23400_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22919__A2 _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21139__B _21139_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23067_ _23047_/X _23050_/X _23054_/Y _23066_/X VGND VGND VPWR VPWR HRDATA[23] sky130_fd_sc_hd__a211o_4
X_20279_ _20275_/Y _20278_/X _19975_/X _20278_/X VGND VGND VPWR VPWR _23427_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12332__A2 _24816_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22018_ _22025_/A _22016_/X _22018_/C VGND VGND VPWR VPWR _22018_/X sky130_fd_sc_hd__and3_4
XFILLER_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15806__B1 _11767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23981__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14840_ _23987_/D _14839_/Y _25184_/Q _23987_/D VGND VGND VPWR VPWR _14840_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21155__A _15336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14771_ _16173_/B _14762_/X _14781_/B VGND VGND VPWR VPWR _14771_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15821__A3 _15745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25134__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11983_ _11654_/B _11976_/X VGND VGND VPWR VPWR _11987_/A sky130_fd_sc_hd__and2_4
XFILLER_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23073__C _22812_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23969_ _24942_/CLK _20608_/Y HRESETn VGND VGND VPWR VPWR _23969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22552__B1 _12305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13722_ _13686_/X _13720_/Y _13721_/X _13714_/X _25274_/Q VGND VGND VPWR VPWR _25274_/D
+ sky130_fd_sc_hd__a32o_4
X_16510_ _16510_/A VGND VGND VPWR VPWR _16510_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17490_ _17480_/Y _17481_/X _17482_/X _17489_/X VGND VGND VPWR VPWR _17491_/A sky130_fd_sc_hd__o22a_4
XFILLER_44_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13653_ _13653_/A _13653_/B VGND VGND VPWR VPWR _13654_/A sky130_fd_sc_hd__and2_4
X_16441_ HWDATA[2] VGND VGND VPWR VPWR _16442_/A sky130_fd_sc_hd__buf_2
XFILLER_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12604_ _12604_/A VGND VGND VPWR VPWR _12665_/A sky130_fd_sc_hd__inv_2
XFILLER_38_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ _16371_/X VGND VGND VPWR VPWR _16728_/B sky130_fd_sc_hd__buf_2
X_19160_ _19153_/Y VGND VGND VPWR VPWR _19160_/X sky130_fd_sc_hd__buf_2
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ _25070_/Q VGND VGND VPWR VPWR _14560_/B sky130_fd_sc_hd__inv_2
XFILLER_125_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15323_ _15309_/C _15320_/X VGND VGND VPWR VPWR _15323_/X sky130_fd_sc_hd__or2_4
X_18111_ _18175_/A _18976_/A VGND VGND VPWR VPWR _18112_/C sky130_fd_sc_hd__or2_4
XFILLER_12_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12535_ _25396_/Q VGND VGND VPWR VPWR _12707_/A sky130_fd_sc_hd__inv_2
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19091_ _19098_/A VGND VGND VPWR VPWR _19091_/X sky130_fd_sc_hd__buf_2
XFILLER_9_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12943__C _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15254_ _14886_/X _15252_/A VGND VGND VPWR VPWR _15254_/X sky130_fd_sc_hd__or2_4
X_18042_ _18080_/A _23874_/Q VGND VGND VPWR VPWR _18042_/X sky130_fd_sc_hd__or2_4
X_12466_ _12465_/X VGND VGND VPWR VPWR _25432_/D sky130_fd_sc_hd__inv_2
XANTENNA__24087__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14205_ _14205_/A VGND VGND VPWR VPWR _14205_/Y sky130_fd_sc_hd__inv_2
X_15185_ _15185_/A VGND VGND VPWR VPWR _15185_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17808__A _17759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24016__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12397_ _12385_/B _12397_/B VGND VGND VPWR VPWR _12398_/A sky130_fd_sc_hd__or2_4
XANTENNA__16712__A _16645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16298__B1 _16297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14136_ _14108_/X VGND VGND VPWR VPWR _14136_/X sky130_fd_sc_hd__buf_2
X_19993_ _19990_/Y _19991_/X _19992_/X _19991_/X VGND VGND VPWR VPWR _23535_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18853__A1_N _16508_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11856__A HWDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14067_ _14001_/D _14065_/X _14057_/X _13999_/X _14066_/X VGND VGND VPWR VPWR _25228_/D
+ sky130_fd_sc_hd__a32o_4
X_18944_ _18944_/A VGND VGND VPWR VPWR _18944_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15328__A _15310_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19236__B1 _19212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13018_ _13012_/A _13017_/X _13010_/A _13013_/Y VGND VGND VPWR VPWR _13019_/A sky130_fd_sc_hd__a211o_4
XFILLER_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18875_ _18875_/A _18875_/B VGND VGND VPWR VPWR _20566_/B sky130_fd_sc_hd__or2_4
XFILLER_121_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17826_ _17826_/A _17826_/B VGND VGND VPWR VPWR _17827_/C sky130_fd_sc_hd__or2_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16470__B1 _16384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13790__B _21027_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21065__A _21065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17757_ _24261_/Q VGND VGND VPWR VPWR _17758_/D sky130_fd_sc_hd__inv_2
XFILLER_78_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14969_ _14969_/A VGND VGND VPWR VPWR _14969_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_13_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__21346__B2 _12096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16708_ _16706_/Y _16707_/X _16528_/X _16707_/X VGND VGND VPWR VPWR _16708_/X sky130_fd_sc_hd__a2bb2o_4
X_17688_ _17578_/C _17695_/A VGND VGND VPWR VPWR _17688_/X sky130_fd_sc_hd__or2_4
XFILLER_39_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16222__B1 _15964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19427_ _19422_/Y _19425_/X _19426_/X _19425_/X VGND VGND VPWR VPWR _23732_/D sky130_fd_sc_hd__a2bb2o_4
X_16639_ _16630_/A _16638_/X _16634_/X VGND VGND VPWR VPWR _24498_/D sky130_fd_sc_hd__o21a_4
XFILLER_126_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24857__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19358_ _17967_/B VGND VGND VPWR VPWR _19358_/Y sky130_fd_sc_hd__inv_2
X_18309_ _21478_/A VGND VGND VPWR VPWR _21658_/A sky130_fd_sc_hd__buf_2
X_19289_ _19284_/Y _19288_/X _19155_/X _19288_/X VGND VGND VPWR VPWR _23780_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21320_ _23170_/A _21320_/B _21320_/C VGND VGND VPWR VPWR _21320_/X sky130_fd_sc_hd__and3_4
XFILLER_15_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13311__A _13227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_137_0_HCLK clkbuf_7_68_0_HCLK/X VGND VGND VPWR VPWR _23660_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21251_ _21247_/X _21250_/X _21233_/X VGND VGND VPWR VPWR _21251_/X sky130_fd_sc_hd__o21a_4
XFILLER_128_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20202_ _23455_/Q VGND VGND VPWR VPWR _20202_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21182_ _21173_/A _20294_/Y VGND VGND VPWR VPWR _21182_/X sky130_fd_sc_hd__or2_4
XFILLER_85_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20133_ _20140_/A VGND VGND VPWR VPWR _20133_/X sky130_fd_sc_hd__buf_2
XANTENNA__23023__A1 _12259_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20064_ _20065_/A VGND VGND VPWR VPWR _20064_/X sky130_fd_sc_hd__buf_2
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24941_ _24148_/CLK _24941_/D HRESETn VGND VGND VPWR VPWR _24941_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21585__A1 _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24872_ _24865_/CLK _24872_/D HRESETn VGND VGND VPWR VPWR _24872_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23823_ _25264_/CLK _23823_/D VGND VGND VPWR VPWR _19166_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_66_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16069__A _24706_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23754_ _23772_/CLK _19362_/X VGND VGND VPWR VPWR _18024_/B sky130_fd_sc_hd__dfxtp_4
X_20966_ _12155_/X _20965_/B VGND VGND VPWR VPWR _20966_/X sky130_fd_sc_hd__and2_4
XANTENNA__16213__B1 _15955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15016__B2 _24434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22705_ _22705_/A _22702_/X _22704_/X VGND VGND VPWR VPWR _22705_/X sky130_fd_sc_hd__and3_4
XFILLER_41_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23685_ _23689_/CLK _23685_/D VGND VGND VPWR VPWR _23685_/Q sky130_fd_sc_hd__dfxtp_4
X_20897_ _24046_/Q _24047_/Q _20889_/A _20889_/B VGND VGND VPWR VPWR _20897_/X sky130_fd_sc_hd__or4_4
XANTENNA__24598__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15701__A _15642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25424_ _25425_/CLK _12497_/Y HRESETn VGND VGND VPWR VPWR _25424_/Q sky130_fd_sc_hd__dfrtp_4
X_22636_ _21580_/A _22636_/B VGND VGND VPWR VPWR _22636_/Y sky130_fd_sc_hd__nor2_4
XFILLER_41_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24527__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25355_ _25330_/CLK _12979_/X HRESETn VGND VGND VPWR VPWR _25355_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_33_0_HCLK clkbuf_7_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_67_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22567_ _12944_/C _22565_/X _22566_/X VGND VGND VPWR VPWR _22567_/X sky130_fd_sc_hd__o21a_4
XFILLER_16_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12250__B2 _24750_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12320_ _25346_/Q VGND VGND VPWR VPWR _13030_/A sky130_fd_sc_hd__inv_2
X_24306_ _24305_/CLK _24306_/D HRESETn VGND VGND VPWR VPWR _24306_/Q sky130_fd_sc_hd__dfrtp_4
X_21518_ _21525_/A VGND VGND VPWR VPWR _21519_/B sky130_fd_sc_hd__buf_2
Xclkbuf_7_96_0_HCLK clkbuf_6_48_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_96_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24180__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25286_ _24026_/CLK _25286_/D HRESETn VGND VGND VPWR VPWR _25286_/Q sky130_fd_sc_hd__dfrtp_4
X_22498_ _15668_/X _22498_/B VGND VGND VPWR VPWR _22498_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22534__A _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12251_ _12243_/X _12245_/X _12251_/C _12250_/X VGND VGND VPWR VPWR _12251_/X sky130_fd_sc_hd__or4_4
XANTENNA__18269__A1 _13795_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24237_ _23516_/CLK _24237_/D HRESETn VGND VGND VPWR VPWR _13541_/B sky130_fd_sc_hd__dfrtp_4
X_21449_ _21449_/A _19509_/Y VGND VGND VPWR VPWR _21449_/X sky130_fd_sc_hd__or2_4
XFILLER_68_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12553__A2 _12552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12182_ _25447_/Q VGND VGND VPWR VPWR _12291_/A sky130_fd_sc_hd__inv_2
X_24168_ _24502_/CLK _18517_/X HRESETn VGND VGND VPWR VPWR _24168_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23119_ _22783_/A VGND VGND VPWR VPWR _23119_/X sky130_fd_sc_hd__buf_2
XANTENNA__25386__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_16990_ _16990_/A _16971_/X _16990_/C _16990_/D VGND VGND VPWR VPWR _16990_/X sky130_fd_sc_hd__or4_4
XANTENNA__23014__B2 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24099_ _23933_/CLK _20964_/X HRESETn VGND VGND VPWR VPWR _12128_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_62_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15941_ _12217_/Y _15939_/X _15940_/X _15939_/X VGND VGND VPWR VPWR _24764_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23365__A _21008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25315__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21576__A1 _16618_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18660_ _18660_/A _18655_/X _18660_/C _18660_/D VGND VGND VPWR VPWR _18667_/C sky130_fd_sc_hd__or4_4
X_15872_ _15868_/X VGND VGND VPWR VPWR _15872_/X sky130_fd_sc_hd__buf_2
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17611_ _17611_/A _17611_/B _17543_/Y _17569_/X VGND VGND VPWR VPWR _17618_/A sky130_fd_sc_hd__or4_4
X_14823_ _14880_/B _14810_/A VGND VGND VPWR VPWR _14824_/A sky130_fd_sc_hd__and2_4
XFILLER_40_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18591_ _18588_/B _18591_/B _18582_/C VGND VGND VPWR VPWR _18591_/X sky130_fd_sc_hd__and3_4
XANTENNA__21328__A1 _16620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17542_ _11759_/Y _24304_/Q _25527_/Q _17541_/Y VGND VGND VPWR VPWR _17545_/C sky130_fd_sc_hd__a2bb2o_4
X_11966_ _11961_/A _11967_/D _11965_/X VGND VGND VPWR VPWR _11966_/Y sky130_fd_sc_hd__a21oi_4
X_14754_ _21612_/A _14752_/X _14753_/Y VGND VGND VPWR VPWR _14754_/X sky130_fd_sc_hd__o21a_4
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13705_ _13693_/A _13693_/B VGND VGND VPWR VPWR _13705_/X sky130_fd_sc_hd__or2_4
X_14685_ _14677_/X _14750_/A _14746_/A VGND VGND VPWR VPWR _14697_/B sky130_fd_sc_hd__o21a_4
X_17473_ _17472_/A _17472_/B _17471_/Y _17472_/Y VGND VGND VPWR VPWR _17473_/X sky130_fd_sc_hd__a211o_4
X_11897_ _11896_/X _11887_/X VGND VGND VPWR VPWR _11897_/Y sky130_fd_sc_hd__nor2_4
XFILLER_32_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24950__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16707__A _16645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19212_ _16442_/A VGND VGND VPWR VPWR _19212_/X sky130_fd_sc_hd__buf_2
X_13636_ _13635_/X VGND VGND VPWR VPWR _13637_/A sky130_fd_sc_hd__buf_2
X_16424_ _16423_/Y _16419_/X _16238_/X _16419_/X VGND VGND VPWR VPWR _24579_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22828__B2 _22827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24268__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19143_ _23831_/Q VGND VGND VPWR VPWR _19143_/Y sky130_fd_sc_hd__inv_2
X_13567_ _13565_/A _13566_/A _13565_/Y _14561_/A VGND VGND VPWR VPWR _13567_/X sky130_fd_sc_hd__o22a_4
X_16355_ _16355_/A VGND VGND VPWR VPWR _16355_/X sky130_fd_sc_hd__buf_2
XFILLER_34_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12518_ _12517_/Y _24867_/Q _12517_/Y _24867_/Q VGND VGND VPWR VPWR _12518_/X sky130_fd_sc_hd__a2bb2o_4
X_15306_ _15336_/D _15336_/B VGND VGND VPWR VPWR _15306_/X sky130_fd_sc_hd__or2_4
XFILLER_118_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16286_ _16284_/Y _16282_/X _16285_/X _16282_/X VGND VGND VPWR VPWR _24629_/D sky130_fd_sc_hd__a2bb2o_4
X_19074_ _19073_/Y _19068_/X _18977_/X _19068_/X VGND VGND VPWR VPWR _19074_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13498_ _13497_/Y VGND VGND VPWR VPWR _13498_/X sky130_fd_sc_hd__buf_2
XFILLER_117_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22444__A _22444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17180__B2 _17242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18025_ _17975_/A VGND VGND VPWR VPWR _18133_/A sky130_fd_sc_hd__buf_2
XFILLER_51_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12449_ _12429_/X _12445_/B _12449_/C VGND VGND VPWR VPWR _12449_/X sky130_fd_sc_hd__and3_4
X_15237_ _15236_/X VGND VGND VPWR VPWR _25009_/D sky130_fd_sc_hd__inv_2
XFILLER_12_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19457__B1 _19389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12970__A _12976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23259__B _23256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23253__B2 _22827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16442__A _16442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15168_ _25026_/Q _15167_/Y VGND VGND VPWR VPWR _15168_/X sky130_fd_sc_hd__or2_4
XFILLER_99_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11752__B1 _11749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14119_ _14119_/A _14118_/Y _14119_/C VGND VGND VPWR VPWR _14120_/B sky130_fd_sc_hd__and3_4
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19209__B1 _19117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15099_ _24575_/Q VGND VGND VPWR VPWR _15099_/Y sky130_fd_sc_hd__inv_2
X_19976_ _22348_/B _19974_/X _19975_/X _19974_/X VGND VGND VPWR VPWR _23540_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16691__B1 _15750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18927_ _18927_/A VGND VGND VPWR VPWR _18927_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25056__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18858_ _16485_/A _18749_/A _24561_/Q _18696_/A VGND VGND VPWR VPWR _18858_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16443__B1 _16442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17809_ _17756_/A _17755_/Y _17830_/B VGND VGND VPWR VPWR _17818_/D sky130_fd_sc_hd__or3_4
XFILLER_83_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18789_ _18789_/A _18788_/Y VGND VGND VPWR VPWR _18791_/B sky130_fd_sc_hd__or2_4
X_20820_ _20819_/X VGND VGND VPWR VPWR _24029_/D sky130_fd_sc_hd__inv_2
XFILLER_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13306__A _13454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12210__A _22400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21523__A _15784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20751_ _20749_/Y _20745_/Y _20750_/X VGND VGND VPWR VPWR _20751_/X sky130_fd_sc_hd__o21a_4
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24691__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23470_ _24089_/CLK _20164_/X VGND VGND VPWR VPWR _23470_/Q sky130_fd_sc_hd__dfxtp_4
X_20682_ _20681_/X VGND VGND VPWR VPWR _23997_/D sky130_fd_sc_hd__inv_2
XANTENNA__24620__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22421_ _22879_/A VGND VGND VPWR VPWR _22421_/X sky130_fd_sc_hd__buf_2
XFILLER_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22295__A2 _22590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25140_ _24943_/CLK _14385_/X HRESETn VGND VGND VPWR VPWR _25140_/Q sky130_fd_sc_hd__dfrtp_4
X_22352_ _17728_/A _22331_/Y _22338_/Y _22345_/Y _22351_/Y VGND VGND VPWR VPWR _22352_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_137_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22354__A _22055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21303_ _22419_/A VGND VGND VPWR VPWR _21303_/X sky130_fd_sc_hd__buf_2
XANTENNA__15182__B1 _15174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17448__A _11710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19382__A2_N _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23244__A1 _24531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25071_ _25070_/CLK _14611_/X HRESETn VGND VGND VPWR VPWR _14610_/A sky130_fd_sc_hd__dfrtp_4
X_22283_ _21741_/A _22283_/B VGND VGND VPWR VPWR _22283_/Y sky130_fd_sc_hd__nor2_4
XFILLER_117_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19448__B1 _19426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16352__A _16352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24022_ _24055_/CLK _24022_/D HRESETn VGND VGND VPWR VPWR _13136_/A sky130_fd_sc_hd__dfrtp_4
X_21234_ _21226_/X _21232_/X _21233_/X VGND VGND VPWR VPWR _21244_/B sky130_fd_sc_hd__o21a_4
XFILLER_116_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21165_ _24200_/Q _21163_/X _21164_/X VGND VGND VPWR VPWR _21165_/X sky130_fd_sc_hd__and3_4
XANTENNA__16277__A3 _16270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22801__B _22801_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20116_ _21756_/B _20111_/X _20092_/X _20111_/X VGND VGND VPWR VPWR _20116_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21096_ _15992_/B VGND VGND VPWR VPWR _22419_/A sky130_fd_sc_hd__buf_2
XFILLER_115_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20047_ _20047_/A VGND VGND VPWR VPWR _20047_/Y sky130_fd_sc_hd__inv_2
X_24924_ _24926_/CLK _15518_/X HRESETn VGND VGND VPWR VPWR _11728_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_85_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16434__B1 _16061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24855_ _24865_/CLK _24855_/D HRESETn VGND VGND VPWR VPWR _24855_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24779__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20781__A2 _20676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11820_ _25517_/Q VGND VGND VPWR VPWR _11820_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13216__A _13454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23806_ _23805_/CLK _23806_/D VGND VGND VPWR VPWR _18190_/B sky130_fd_sc_hd__dfxtp_4
X_24786_ _24800_/CLK _24786_/D HRESETn VGND VGND VPWR VPWR _22708_/A sky130_fd_sc_hd__dfrtp_4
X_21998_ _20385_/Y _21995_/Y _22384_/A _21997_/Y VGND VGND VPWR VPWR _21998_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24708__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21433__A _21433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11777_/A VGND VGND VPWR VPWR _11751_/X sky130_fd_sc_hd__buf_2
XPHY_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23737_ _23718_/CLK _23737_/D VGND VGND VPWR VPWR _23737_/Q sky130_fd_sc_hd__dfxtp_4
X_20949_ _20818_/X _20948_/X _24496_/Q _20864_/X VGND VGND VPWR VPWR _24059_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16527__A _24539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _14470_/A VGND VGND VPWR VPWR _14470_/X sky130_fd_sc_hd__buf_2
XPHY_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11682_/A VGND VGND VPWR VPWR _11682_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24361__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23668_ _23580_/CLK _23668_/D VGND VGND VPWR VPWR _23668_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13421_/A _13419_/X _13421_/C VGND VGND VPWR VPWR _13421_/X sky130_fd_sc_hd__and3_4
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25407_ _25020_/CLK _25407_/D HRESETn VGND VGND VPWR VPWR _25407_/Q sky130_fd_sc_hd__dfrtp_4
X_22619_ _22619_/A _22522_/B VGND VGND VPWR VPWR _22619_/X sky130_fd_sc_hd__or2_4
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23599_ _23598_/CLK _19816_/X VGND VGND VPWR VPWR _23599_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16140_ _22556_/A VGND VGND VPWR VPWR _16140_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13352_ _13316_/A _19673_/A VGND VGND VPWR VPWR _13354_/B sky130_fd_sc_hd__or2_4
XANTENNA__21494__B1 _21493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25338_ _24852_/CLK _25338_/D HRESETn VGND VGND VPWR VPWR _12302_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22264__A _21275_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12303_ _12303_/A VGND VGND VPWR VPWR _13057_/A sky130_fd_sc_hd__buf_2
X_16071_ _24705_/Q VGND VGND VPWR VPWR _16071_/Y sky130_fd_sc_hd__inv_2
X_13283_ _13320_/A _23658_/Q VGND VGND VPWR VPWR _13283_/X sky130_fd_sc_hd__or2_4
XANTENNA__19439__B1 _19370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17358__A _17350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25269_ _24214_/CLK _25269_/D HRESETn VGND VGND VPWR VPWR _11682_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_120_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15022_ _15022_/A _15002_/X _15012_/X _15021_/X VGND VGND VPWR VPWR _15022_/X sky130_fd_sc_hd__or4_4
Xclkbuf_8_120_0_HCLK clkbuf_7_60_0_HCLK/X VGND VGND VPWR VPWR _24654_/CLK sky130_fd_sc_hd__clkbuf_1
X_12234_ _25432_/Q VGND VGND VPWR VPWR _12235_/A sky130_fd_sc_hd__inv_2
Xclkbuf_8_183_0_HCLK clkbuf_7_91_0_HCLK/X VGND VGND VPWR VPWR _24759_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19830_ _19828_/Y _19824_/X _19783_/X _19829_/X VGND VGND VPWR VPWR _23594_/D sky130_fd_sc_hd__a2bb2o_4
X_12165_ _24094_/Q VGND VGND VPWR VPWR _14325_/A sky130_fd_sc_hd__inv_2
XFILLER_110_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23095__A _21108_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19761_ _23617_/Q VGND VGND VPWR VPWR _19761_/Y sky130_fd_sc_hd__inv_2
X_12096_ _12095_/Y VGND VGND VPWR VPWR _12096_/X sky130_fd_sc_hd__buf_2
X_16973_ _24722_/Q _24379_/Q _16026_/Y _16972_/Y VGND VGND VPWR VPWR _16973_/X sky130_fd_sc_hd__o22a_4
XFILLER_42_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13487__B1 _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18712_ _24142_/Q _18712_/B VGND VGND VPWR VPWR _18714_/B sky130_fd_sc_hd__or2_4
X_15924_ _15646_/X _15835_/X _15845_/X _21005_/B _15923_/X VGND VGND VPWR VPWR _15924_/X
+ sky130_fd_sc_hd__a32o_4
X_19692_ _13317_/B VGND VGND VPWR VPWR _19692_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18643_ _16592_/Y _18686_/A _16592_/Y _18686_/A VGND VGND VPWR VPWR _18643_/X sky130_fd_sc_hd__a2bb2o_4
X_15855_ _15854_/X VGND VGND VPWR VPWR _15894_/A sky130_fd_sc_hd__buf_2
XFILLER_76_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14806_ _14819_/C _14806_/B _14820_/A VGND VGND VPWR VPWR _14807_/C sky130_fd_sc_hd__and3_4
XFILLER_92_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18574_ _18555_/A _18574_/B _18573_/Y VGND VGND VPWR VPWR _24153_/D sky130_fd_sc_hd__and3_4
X_15786_ _15925_/B VGND VGND VPWR VPWR _15819_/A sky130_fd_sc_hd__inv_2
XFILLER_79_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24449__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12998_ _13028_/D _13043_/B VGND VGND VPWR VPWR _12999_/D sky130_fd_sc_hd__or2_4
XANTENNA__22439__A _21306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17525_ _24295_/Q VGND VGND VPWR VPWR _17525_/Y sky130_fd_sc_hd__inv_2
X_14737_ _14733_/Y _14736_/Y _14732_/X _14736_/A VGND VGND VPWR VPWR _14737_/X sky130_fd_sc_hd__o22a_4
X_11949_ _11946_/Y _11947_/X _11948_/X _11947_/X VGND VGND VPWR VPWR _25492_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12247__A1_N _12286_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16548__A1_N _16547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17456_ _17456_/A VGND VGND VPWR VPWR _17456_/Y sky130_fd_sc_hd__inv_2
X_14668_ _14659_/A _14667_/X _19014_/B _13633_/B VGND VGND VPWR VPWR _14668_/X sky130_fd_sc_hd__o22a_4
X_16407_ _15096_/Y _16400_/X _16405_/X _16406_/X VGND VGND VPWR VPWR _24586_/D sky130_fd_sc_hd__a2bb2o_4
X_13619_ _13617_/Y _13618_/Y VGND VGND VPWR VPWR _13619_/X sky130_fd_sc_hd__or2_4
X_17387_ _17387_/A VGND VGND VPWR VPWR _17387_/X sky130_fd_sc_hd__buf_2
XANTENNA__24031__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14599_ _14586_/A VGND VGND VPWR VPWR _14599_/X sky130_fd_sc_hd__buf_2
X_19126_ _19126_/A VGND VGND VPWR VPWR _19126_/Y sky130_fd_sc_hd__inv_2
X_16338_ _16336_/Y _16337_/X _16242_/X _16337_/X VGND VGND VPWR VPWR _24610_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12800__A1_N _12799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11973__B1 _11958_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19057_ _19054_/Y _19052_/X _19056_/X _19052_/X VGND VGND VPWR VPWR _23862_/D sky130_fd_sc_hd__a2bb2o_4
X_16269_ _16268_/Y _16187_/A _15480_/X _16187_/A VGND VGND VPWR VPWR _16269_/X sky130_fd_sc_hd__a2bb2o_4
X_18008_ _18088_/A VGND VGND VPWR VPWR _18150_/A sky130_fd_sc_hd__buf_2
XANTENNA__25237__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18653__B2 _18608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21518__A _21525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19959_ _23545_/Q VGND VGND VPWR VPWR _21929_/B sky130_fd_sc_hd__inv_2
XANTENNA__13478__B1 _11833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22970_ _22897_/A _22970_/B VGND VGND VPWR VPWR _22979_/C sky130_fd_sc_hd__and2_4
XFILLER_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12150__B1 _12104_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21921_ _21917_/X _21921_/B _21921_/C VGND VGND VPWR VPWR _21921_/X sky130_fd_sc_hd__and3_4
XFILLER_132_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24872__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24640_ _24162_/CLK _16255_/X HRESETn VGND VGND VPWR VPWR _22154_/A sky130_fd_sc_hd__dfrtp_4
X_21852_ _21852_/A _22695_/B _22695_/C VGND VGND VPWR VPWR _21852_/X sky130_fd_sc_hd__and3_4
XFILLER_58_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24801__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20803_ _20804_/A VGND VGND VPWR VPWR _20803_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24571_ _24572_/CLK _16438_/X HRESETn VGND VGND VPWR VPWR _24571_/Q sky130_fd_sc_hd__dfrtp_4
X_21783_ _21782_/X VGND VGND VPWR VPWR _21783_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24119__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23522_ _23714_/CLK _23522_/D VGND VGND VPWR VPWR _20028_/A sky130_fd_sc_hd__dfxtp_4
X_20734_ _13133_/A VGND VGND VPWR VPWR _20734_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12205__A1 _12202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23453_ _23453_/CLK _20208_/X VGND VGND VPWR VPWR _23453_/Q sky130_fd_sc_hd__dfxtp_4
X_20665_ _20488_/B _20665_/B _20665_/C VGND VGND VPWR VPWR _20665_/X sky130_fd_sc_hd__and3_4
XANTENNA__19658__A _15845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12205__B2 _12204_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22404_ _21064_/X _22401_/X _22270_/X _22403_/X VGND VGND VPWR VPWR _22405_/B sky130_fd_sc_hd__a22oi_4
XFILLER_52_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23384_ _23384_/CLK _23384_/D VGND VGND VPWR VPWR _23384_/Q sky130_fd_sc_hd__dfxtp_4
X_20596_ _20596_/A _20443_/B VGND VGND VPWR VPWR _20596_/X sky130_fd_sc_hd__or2_4
X_25123_ _25113_/CLK _25123_/D HRESETn VGND VGND VPWR VPWR _25123_/Q sky130_fd_sc_hd__dfstp_4
X_22335_ _21929_/A _19949_/Y VGND VGND VPWR VPWR _22337_/B sky130_fd_sc_hd__or2_4
XFILLER_109_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23217__B2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25054_ _25054_/CLK _14739_/X HRESETn VGND VGND VPWR VPWR _25054_/Q sky130_fd_sc_hd__dfrtp_4
X_22266_ _22590_/B VGND VGND VPWR VPWR _22266_/X sky130_fd_sc_hd__buf_2
XFILLER_133_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21779__A1 _21636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22812__A _24551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21779__B2 _18261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24005_ _24035_/CLK _20716_/Y HRESETn VGND VGND VPWR VPWR _20712_/A sky130_fd_sc_hd__dfrtp_4
X_21217_ _21018_/A VGND VGND VPWR VPWR _21323_/A sky130_fd_sc_hd__buf_2
XFILLER_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22197_ _22200_/A _22197_/B VGND VGND VPWR VPWR _22197_/X sky130_fd_sc_hd__or2_4
X_21148_ _17438_/Y _21116_/Y _14190_/B _21147_/X VGND VGND VPWR VPWR _21148_/X sky130_fd_sc_hd__a211o_4
XFILLER_28_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13970_ _13970_/A _13944_/Y _13970_/C _13962_/Y VGND VGND VPWR VPWR _13971_/A sky130_fd_sc_hd__or4_4
X_21079_ _21005_/A _21038_/B VGND VGND VPWR VPWR _21079_/X sky130_fd_sc_hd__and2_4
XFILLER_101_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16407__B1 _16405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12921_ _12936_/A _12917_/B _12920_/X VGND VGND VPWR VPWR _25372_/D sky130_fd_sc_hd__and3_4
XANTENNA__22743__A3 _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24907_ _24055_/CLK _15571_/X HRESETn VGND VGND VPWR VPWR _15570_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_98_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20986__B _14196_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17080__B1 _17056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15640_ _12049_/A _15640_/B _15700_/C _15549_/X VGND VGND VPWR VPWR _15641_/A sky130_fd_sc_hd__or4_4
XFILLER_34_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12852_ _12847_/X _12852_/B VGND VGND VPWR VPWR _12852_/X sky130_fd_sc_hd__or2_4
X_24838_ _24830_/CLK _15794_/X HRESETn VGND VGND VPWR VPWR _24838_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24542__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23153__B1 _25533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18456__B _18503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11803_ HWDATA[14] VGND VGND VPWR VPWR _11803_/X sky130_fd_sc_hd__buf_2
X_12783_ _12871_/A _24801_/Q _12864_/A _12782_/Y VGND VGND VPWR VPWR _12783_/X sky130_fd_sc_hd__o22a_4
X_15571_ _15570_/Y _15568_/X _11757_/X _15568_/X VGND VGND VPWR VPWR _15571_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ _24806_/CLK _15924_/X HRESETn VGND VGND VPWR VPWR _21005_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__22900__B1 _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17220_/Y _17309_/X VGND VGND VPWR VPWR _17311_/A sky130_fd_sc_hd__or2_4
XFILLER_15_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11734_ _11734_/A VGND VGND VPWR VPWR _21314_/A sky130_fd_sc_hd__inv_2
X_14522_ _25094_/Q _14511_/X _21841_/A _14513_/X VGND VGND VPWR VPWR _14522_/X sky130_fd_sc_hd__o22a_4
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18290_ _24198_/Q _19492_/B _17700_/X VGND VGND VPWR VPWR _18300_/A sky130_fd_sc_hd__a21o_4
XPHY_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _24332_/Q VGND VGND VPWR VPWR _17348_/A sky130_fd_sc_hd__inv_2
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11663_/Y _24219_/Q _13676_/A _11664_/Y VGND VGND VPWR VPWR _11666_/D sky130_fd_sc_hd__a2bb2o_4
X_14453_ _15851_/B _14475_/B VGND VGND VPWR VPWR _14453_/Y sky130_fd_sc_hd__nor2_4
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22706__B _21220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _13303_/A _13404_/B VGND VGND VPWR VPWR _13404_/X sky130_fd_sc_hd__or2_4
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ _14384_/A VGND VGND VPWR VPWR _14384_/X sky130_fd_sc_hd__buf_2
X_17172_ _17172_/A _17172_/B _17170_/X _17171_/X VGND VGND VPWR VPWR _17202_/A sky130_fd_sc_hd__or4_4
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20507__A _14205_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13335_ _13198_/X _13334_/X _25317_/Q _13258_/X VGND VGND VPWR VPWR _25317_/D sky130_fd_sc_hd__o22a_4
X_16123_ _16122_/Y _16118_/X _15964_/X _16118_/X VGND VGND VPWR VPWR _24685_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17088__A _17384_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13266_ _13373_/A _13266_/B VGND VGND VPWR VPWR _13267_/C sky130_fd_sc_hd__or2_4
X_16054_ _24711_/Q VGND VGND VPWR VPWR _16054_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25330__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15541__A2_N _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22100__A2_N _21548_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12217_ _24764_/Q VGND VGND VPWR VPWR _12217_/Y sky130_fd_sc_hd__inv_2
X_15005_ _15005_/A VGND VGND VPWR VPWR _15005_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13197_ _13176_/X _13193_/X _13195_/X _25320_/Q _13196_/Y VGND VGND VPWR VPWR _25320_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22431__A2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19832__B1 _19787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19813_ _19812_/Y _19808_/X _19740_/X _19808_/X VGND VGND VPWR VPWR _19813_/X sky130_fd_sc_hd__a2bb2o_4
X_12148_ _12148_/A VGND VGND VPWR VPWR _12148_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21338__A _14220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19744_ _19742_/Y _19743_/X _19721_/X _19743_/X VGND VGND VPWR VPWR _19744_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15336__A _15336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12079_ _12073_/Y VGND VGND VPWR VPWR _12079_/X sky130_fd_sc_hd__buf_2
X_16956_ _24700_/Q VGND VGND VPWR VPWR _16956_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17254__C _17254_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18399__B1 _16199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15907_ _15705_/X _15894_/X _15768_/X _24775_/Q _15864_/A VGND VGND VPWR VPWR _15907_/X
+ sky130_fd_sc_hd__a32o_4
X_19675_ _23647_/Q VGND VGND VPWR VPWR _19675_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16887_ _19841_/A VGND VGND VPWR VPWR _16887_/Y sky130_fd_sc_hd__inv_2
X_18626_ _24132_/Q VGND VGND VPWR VPWR _18626_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15838_ _15824_/X _15835_/X _15768_/X _24810_/Q _15793_/A VGND VGND VPWR VPWR _15838_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24283__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21073__A _24735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18557_ _18556_/X VGND VGND VPWR VPWR _24157_/D sky130_fd_sc_hd__inv_2
X_15769_ _15749_/X _15765_/X _15768_/X _24845_/Q _15711_/A VGND VGND VPWR VPWR _15769_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_17_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17508_ _24286_/Q VGND VGND VPWR VPWR _17676_/A sky130_fd_sc_hd__inv_2
XFILLER_33_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18488_ _18482_/A _18482_/B _18483_/B _18487_/X VGND VGND VPWR VPWR _18489_/A sky130_fd_sc_hd__a211o_4
XFILLER_36_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17439_ _12095_/Y _13789_/D _15662_/B VGND VGND VPWR VPWR _17439_/X sky130_fd_sc_hd__or3_4
XANTENNA__25489__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20450_ _23993_/Q _20512_/B _20443_/X _20449_/Y VGND VGND VPWR VPWR _20450_/X sky130_fd_sc_hd__a211o_4
XFILLER_20_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25418__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19109_ _13206_/B VGND VGND VPWR VPWR _19109_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20381_ _20380_/X VGND VGND VPWR VPWR _20381_/X sky130_fd_sc_hd__buf_2
X_22120_ _21306_/X VGND VGND VPWR VPWR _22132_/A sky130_fd_sc_hd__buf_2
XANTENNA__20681__A1 _15638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12124__A1_N _12123_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20681__B2 _20680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25071__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22051_ _22050_/X _19828_/Y VGND VGND VPWR VPWR _22053_/B sky130_fd_sc_hd__or2_4
XANTENNA__25000__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21002_ _24312_/Q _23955_/Q VGND VGND VPWR VPWR _21002_/X sky130_fd_sc_hd__and2_4
XFILLER_138_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_23_0_HCLK clkbuf_8_22_0_HCLK/A VGND VGND VPWR VPWR _25205_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22870__A1_N _17254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15246__A _15246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11774__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_86_0_HCLK clkbuf_8_87_0_HCLK/A VGND VGND VPWR VPWR _24069_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_101_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22953_ _22819_/X _22944_/Y _22948_/Y _22952_/X VGND VGND VPWR VPWR _22961_/C sky130_fd_sc_hd__a211o_4
XFILLER_21_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21904_ _21904_/A _21904_/B VGND VGND VPWR VPWR _21905_/C sky130_fd_sc_hd__or2_4
XFILLER_44_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22884_ _24585_/Q _22884_/B VGND VGND VPWR VPWR _22884_/X sky130_fd_sc_hd__or2_4
X_21835_ _21302_/X _21825_/X _21834_/X VGND VGND VPWR VPWR _21984_/A sky130_fd_sc_hd__a21bo_4
X_24623_ _24355_/CLK _24623_/D HRESETn VGND VGND VPWR VPWR _23073_/A sky130_fd_sc_hd__dfrtp_4
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24554_ _24555_/CLK _24554_/D HRESETn VGND VGND VPWR VPWR _24554_/Q sky130_fd_sc_hd__dfrtp_4
X_21766_ _21624_/A _21766_/B _21766_/C VGND VGND VPWR VPWR _21766_/X sky130_fd_sc_hd__and3_4
XFILLER_19_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14179__A1 _14177_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20717_ _20717_/A VGND VGND VPWR VPWR _20717_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15376__B1 _15318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23505_ _24208_/CLK _23505_/D VGND VGND VPWR VPWR _13312_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24485_ _24447_/CLK _24485_/D HRESETn VGND VGND VPWR VPWR _24485_/Q sky130_fd_sc_hd__dfrtp_4
X_21697_ _24738_/Q _22879_/A VGND VGND VPWR VPWR _21697_/X sky130_fd_sc_hd__or2_4
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18292__A _21192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23935__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23436_ _23434_/CLK _23436_/D VGND VGND VPWR VPWR _23436_/Q sky130_fd_sc_hd__dfxtp_4
X_20648_ _14233_/Y _20628_/X _20619_/A _20647_/X VGND VGND VPWR VPWR _20648_/X sky130_fd_sc_hd__a211o_4
XANTENNA__25159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22110__A1 _21306_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23367_ _23967_/CLK scl_oen_o_S5 VGND VGND VPWR VPWR _23367_/Q sky130_fd_sc_hd__dfxtp_4
X_20579_ _18879_/X _20579_/B _20571_/C VGND VGND VPWR VPWR _20579_/X sky130_fd_sc_hd__and3_4
XANTENNA__22661__A2 _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13120_ _13120_/A _13120_/B _24019_/Q _13120_/D VGND VGND VPWR VPWR _13120_/X sky130_fd_sc_hd__or4_4
X_22318_ _22318_/A VGND VGND VPWR VPWR _22318_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25106_ _25113_/CLK _25106_/D HRESETn VGND VGND VPWR VPWR _14480_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23298_ _23207_/A _23295_/X _23298_/C VGND VGND VPWR VPWR _23299_/D sky130_fd_sc_hd__and3_4
X_13051_ _13050_/X VGND VGND VPWR VPWR _25342_/D sky130_fd_sc_hd__inv_2
X_25037_ _24171_/CLK _14848_/X HRESETn VGND VGND VPWR VPWR _25037_/Q sky130_fd_sc_hd__dfrtp_4
X_22249_ _18293_/B _22249_/B VGND VGND VPWR VPWR _22249_/X sky130_fd_sc_hd__or2_4
XFILLER_65_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12002_ _25298_/Q _12001_/A _12000_/Y _12001_/Y VGND VGND VPWR VPWR _12002_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17355__B _17350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24794__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16810_ _16809_/Y _16807_/X _15725_/X _16807_/X VGND VGND VPWR VPWR _16810_/X sky130_fd_sc_hd__a2bb2o_4
X_17790_ _17790_/A _17790_/B _17790_/C VGND VGND VPWR VPWR _17791_/A sky130_fd_sc_hd__or3_4
XFILLER_59_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24723__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16741_ _24458_/Q VGND VGND VPWR VPWR _16741_/Y sky130_fd_sc_hd__inv_2
X_13953_ _13953_/A _13947_/A _13946_/D VGND VGND VPWR VPWR _13968_/A sky130_fd_sc_hd__or3_4
X_12904_ _12851_/D _12903_/X VGND VGND VPWR VPWR _12905_/B sky130_fd_sc_hd__or2_4
X_19460_ _19458_/Y _19459_/X _19370_/X _19459_/X VGND VGND VPWR VPWR _19460_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16672_ _16670_/Y _16671_/X _16403_/X _16671_/X VGND VGND VPWR VPWR _24486_/D sky130_fd_sc_hd__a2bb2o_4
X_13884_ _14249_/A VGND VGND VPWR VPWR _20467_/A sky130_fd_sc_hd__buf_2
X_18411_ _24152_/Q VGND VGND VPWR VPWR _18411_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16800__B1 _15714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15623_ _15623_/A VGND VGND VPWR VPWR _15623_/X sky130_fd_sc_hd__buf_2
X_12835_ _12829_/X _12831_/X _12832_/X _12835_/D VGND VGND VPWR VPWR _12836_/D sky130_fd_sc_hd__or4_4
X_19391_ _18133_/B VGND VGND VPWR VPWR _19391_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18342_ _17453_/B _18338_/X VGND VGND VPWR VPWR _18345_/A sky130_fd_sc_hd__and2_4
X_15554_ _11734_/A VGND VGND VPWR VPWR _21154_/B sky130_fd_sc_hd__buf_2
X_12766_ _25373_/Q _22857_/A _12764_/Y _12765_/Y VGND VGND VPWR VPWR _12766_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17356__A1 _17350_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14513_/A VGND VGND VPWR VPWR _14505_/X sky130_fd_sc_hd__buf_2
XANTENNA__21621__A _21616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11717_ _12052_/A VGND VGND VPWR VPWR _15549_/A sky130_fd_sc_hd__inv_2
X_18273_ _13784_/D _18237_/A _11867_/A _13695_/A _18272_/X VGND VGND VPWR VPWR _18273_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _12570_/Y _12695_/A VGND VGND VPWR VPWR _12697_/X sky130_fd_sc_hd__or2_4
X_15485_ HTRANS[1] VGND VGND VPWR VPWR _15485_/Y sky130_fd_sc_hd__inv_2
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17224_ _17224_/A _17224_/B _17221_/X _17223_/X VGND VGND VPWR VPWR _17224_/X sky130_fd_sc_hd__or4_4
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _24311_/Q VGND VGND VPWR VPWR _17481_/C sky130_fd_sc_hd__inv_2
X_14436_ _15462_/A _18895_/A VGND VGND VPWR VPWR _14436_/Y sky130_fd_sc_hd__nor2_4
XFILLER_30_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25511__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17155_ _16985_/Y _17159_/B VGND VGND VPWR VPWR _17160_/A sky130_fd_sc_hd__or2_4
XANTENNA__20112__B1 _20085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14367_ _14354_/Y _14366_/X _12083_/A _14360_/X VGND VGND VPWR VPWR _25144_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18856__B2 _18675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24038__CLK _24581_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18930__A _18937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16106_ _16094_/A VGND VGND VPWR VPWR _16106_/X sky130_fd_sc_hd__buf_2
X_13318_ _13386_/A _13318_/B _13318_/C VGND VGND VPWR VPWR _13322_/B sky130_fd_sc_hd__and3_4
XANTENNA__21860__B1 _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14298_ _14291_/A _14301_/B _14297_/Y VGND VGND VPWR VPWR _14298_/X sky130_fd_sc_hd__o21a_4
X_17086_ _17064_/A _17086_/B _17086_/C VGND VGND VPWR VPWR _24383_/D sky130_fd_sc_hd__and3_4
X_16037_ _16037_/A VGND VGND VPWR VPWR _16037_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12568__A2_N _24856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13249_ _13452_/A _23627_/Q VGND VGND VPWR VPWR _13249_/X sky130_fd_sc_hd__or2_4
XFILLER_87_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22404__A2 _22401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16619__B1 _16442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21068__A _21154_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17988_ _17996_/A VGND VGND VPWR VPWR _18211_/A sky130_fd_sc_hd__buf_2
XANTENNA__24464__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12105__B1 _11829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15842__A1 _15824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20058__A1_N _20056_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19727_ _23628_/Q VGND VGND VPWR VPWR _19727_/Y sky130_fd_sc_hd__inv_2
X_16939_ _24273_/Q VGND VGND VPWR VPWR _16939_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19658_ _15845_/A VGND VGND VPWR VPWR _19658_/X sky130_fd_sc_hd__buf_2
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18609_ _16597_/A _18608_/X _16557_/Y _24139_/Q VGND VGND VPWR VPWR _18616_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19589_ _19580_/Y _19588_/X _19426_/X _19588_/X VGND VGND VPWR VPWR _19589_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21620_ _21250_/A VGND VGND VPWR VPWR _21624_/A sky130_fd_sc_hd__buf_2
X_21551_ _21550_/Y _21143_/X _14868_/Y _21352_/X VGND VGND VPWR VPWR _21552_/A sky130_fd_sc_hd__o22a_4
XFILLER_33_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15358__B1 _15318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20502_ _20502_/A VGND VGND VPWR VPWR _20503_/B sky130_fd_sc_hd__inv_2
XFILLER_18_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24270_ _24691_/CLK _17798_/X HRESETn VGND VGND VPWR VPWR _17742_/A sky130_fd_sc_hd__dfrtp_4
X_21482_ _21475_/X _21480_/X _21481_/X VGND VGND VPWR VPWR _21482_/X sky130_fd_sc_hd__o21a_4
XFILLER_21_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25252__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23221_ _23105_/X _23218_/Y _23150_/X _23220_/X VGND VGND VPWR VPWR _23221_/X sky130_fd_sc_hd__a2bb2o_4
X_20433_ _20431_/Y VGND VGND VPWR VPWR _20433_/X sky130_fd_sc_hd__buf_2
X_23152_ _24694_/Q _23310_/B VGND VGND VPWR VPWR _23152_/X sky130_fd_sc_hd__or2_4
X_20364_ _22234_/B _20361_/X _19615_/A _20361_/X VGND VGND VPWR VPWR _23394_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22103_ _15641_/A VGND VGND VPWR VPWR _22103_/X sky130_fd_sc_hd__buf_2
XFILLER_134_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15530__B1 HADDR[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23083_ _24457_/Q _23019_/B _23019_/C VGND VGND VPWR VPWR _23083_/X sky130_fd_sc_hd__and3_4
X_20295_ _20294_/Y _20290_/X _20019_/X _20290_/A VGND VGND VPWR VPWR _23420_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22034_ _21821_/A _21993_/Y _22000_/X _21502_/X _22033_/X VGND VGND VPWR VPWR _22034_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_130_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22159__B2 _21355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24134__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13844__B1 _13800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23985_ _23964_/CLK sda_i_S5 HRESETn VGND VGND VPWR VPWR _23985_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22936_ _24554_/Q _22810_/X _23005_/C VGND VGND VPWR VPWR _22936_/X sky130_fd_sc_hd__and3_4
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22867_ _22769_/X _22862_/Y _22863_/X _22866_/X VGND VGND VPWR VPWR _22867_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13224__A _13233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12620_ _12651_/A _12620_/B _12620_/C _12619_/X VGND VGND VPWR VPWR _12620_/X sky130_fd_sc_hd__or4_4
XFILLER_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24606_ _24606_/CLK _16348_/X HRESETn VGND VGND VPWR VPWR _22402_/A sky130_fd_sc_hd__dfrtp_4
X_21818_ _21636_/X _21817_/X _24211_/Q _21264_/X VGND VGND VPWR VPWR _21818_/X sky130_fd_sc_hd__o22a_4
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22798_ _22798_/A VGND VGND VPWR VPWR _22798_/X sky130_fd_sc_hd__buf_2
XFILLER_12_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21134__A2 _24178_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ _25390_/Q VGND VGND VPWR VPWR _12729_/A sky130_fd_sc_hd__inv_2
X_21749_ _21630_/A _21749_/B VGND VGND VPWR VPWR _21749_/X sky130_fd_sc_hd__or2_4
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24537_ _24545_/CLK _24537_/D HRESETn VGND VGND VPWR VPWR _24537_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _25429_/Q _12481_/Y VGND VGND VPWR VPWR _12482_/X sky130_fd_sc_hd__or2_4
X_15270_ _15267_/A _15267_/B VGND VGND VPWR VPWR _15271_/C sky130_fd_sc_hd__nand2_4
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24468_ _24033_/CLK _24468_/D HRESETn VGND VGND VPWR VPWR _16714_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14221_ _14221_/A VGND VGND VPWR VPWR _14223_/A sky130_fd_sc_hd__buf_2
XFILLER_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23419_ _23394_/CLK _23419_/D VGND VGND VPWR VPWR _23419_/Q sky130_fd_sc_hd__dfxtp_4
X_24399_ _24398_/CLK _24399_/D HRESETn VGND VGND VPWR VPWR _16861_/A sky130_fd_sc_hd__dfrtp_4
X_14152_ _14144_/X _14151_/Y _25205_/Q _14144_/X VGND VGND VPWR VPWR _14152_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16849__B1 _16782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19259__A1_N _21373_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22272__A _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24975__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13103_ _13082_/X _13103_/B _13115_/C VGND VGND VPWR VPWR _25327_/D sky130_fd_sc_hd__and3_4
XANTENNA__14324__A1 _14329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22703__C _21859_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14083_ _13980_/A _14081_/X _14078_/X _13977_/X _14076_/X VGND VGND VPWR VPWR _25220_/D
+ sky130_fd_sc_hd__a32o_4
X_18960_ _18946_/Y VGND VGND VPWR VPWR _18960_/X sky130_fd_sc_hd__buf_2
XFILLER_98_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16270__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24904__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13034_ _13030_/A _13038_/B VGND VGND VPWR VPWR _13034_/Y sky130_fd_sc_hd__nand2_4
X_17911_ _17911_/A VGND VGND VPWR VPWR _17911_/Y sky130_fd_sc_hd__inv_2
X_18891_ _18869_/X _18883_/X _24106_/Q _24107_/Q _18886_/X VGND VGND VPWR VPWR _18891_/X
+ sky130_fd_sc_hd__a32o_4
X_17842_ _17834_/A _17840_/X _17842_/C VGND VGND VPWR VPWR _24258_/D sky130_fd_sc_hd__and3_4
XFILLER_26_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21616__A _21616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17773_ _17765_/C _17772_/X _16955_/X _17768_/B VGND VGND VPWR VPWR _17774_/A sky130_fd_sc_hd__a211o_4
X_14985_ _14940_/X _14984_/X VGND VGND VPWR VPWR _14986_/A sky130_fd_sc_hd__or2_4
XFILLER_47_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18197__A _18010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19512_ _21181_/B _19507_/X _19488_/X _19494_/Y VGND VGND VPWR VPWR _19512_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16724_ _23021_/A VGND VGND VPWR VPWR _22574_/A sky130_fd_sc_hd__buf_2
XFILLER_35_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13936_ _13936_/A VGND VGND VPWR VPWR _13964_/B sky130_fd_sc_hd__inv_2
XFILLER_47_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19443_ _19442_/Y _19438_/X _19420_/X _19431_/A VGND VGND VPWR VPWR _19443_/X sky130_fd_sc_hd__a2bb2o_4
X_16655_ _24492_/Q VGND VGND VPWR VPWR _16655_/Y sky130_fd_sc_hd__inv_2
X_13867_ _13856_/Y VGND VGND VPWR VPWR _13867_/X sky130_fd_sc_hd__buf_2
XANTENNA__18925__A _18937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15606_ _15604_/Y _15600_/X _11809_/X _15605_/X VGND VGND VPWR VPWR _15606_/X sky130_fd_sc_hd__a2bb2o_4
X_12818_ _25359_/Q VGND VGND VPWR VPWR _12819_/A sky130_fd_sc_hd__inv_2
X_19374_ _18196_/B VGND VGND VPWR VPWR _19374_/Y sky130_fd_sc_hd__inv_2
X_16586_ _16585_/Y _16583_/X _16228_/X _16583_/X VGND VGND VPWR VPWR _24517_/D sky130_fd_sc_hd__a2bb2o_4
X_13798_ _23336_/A _13796_/X _13797_/X _13796_/X VGND VGND VPWR VPWR _13798_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22447__A _15668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14260__B1 _13835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18325_ _18325_/A VGND VGND VPWR VPWR _18325_/X sky130_fd_sc_hd__buf_2
X_15537_ _13496_/B _15535_/X HADDR[3] _15535_/X VGND VGND VPWR VPWR _15537_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12749_ _12749_/A VGND VGND VPWR VPWR _12749_/Y sky130_fd_sc_hd__inv_2
X_18256_ _11694_/Y _18249_/X _16852_/X _18233_/A VGND VGND VPWR VPWR _24215_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15468_ _15476_/A VGND VGND VPWR VPWR _15468_/X sky130_fd_sc_hd__buf_2
X_17207_ _24333_/Q VGND VGND VPWR VPWR _17365_/A sky130_fd_sc_hd__inv_2
X_14419_ _14408_/Y VGND VGND VPWR VPWR _14419_/X sky130_fd_sc_hd__buf_2
XANTENNA__22086__B1 _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18187_ _18187_/A _19169_/A VGND VGND VPWR VPWR _18188_/C sky130_fd_sc_hd__or2_4
XANTENNA__15760__B1 _15758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15399_ _15384_/A _15399_/B _15398_/Y VGND VGND VPWR VPWR _24973_/D sky130_fd_sc_hd__and3_4
XFILLER_11_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20636__A1 _14241_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17138_ _17041_/D _17135_/B VGND VGND VPWR VPWR _17138_/Y sky130_fd_sc_hd__nand2_4
XFILLER_85_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17276__A _23246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17069_ _17068_/X VGND VGND VPWR VPWR _24388_/D sky130_fd_sc_hd__inv_2
XANTENNA__15512__B1 HADDR[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24645__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20080_ _22371_/B _20078_/X _20079_/X _20078_/X VGND VGND VPWR VPWR _23500_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21526__A _21526_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13826__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15524__A _15535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23770_ _25503_/CLK _23770_/D VGND VGND VPWR VPWR _19317_/A sky130_fd_sc_hd__dfxtp_4
X_20982_ _20982_/A _20982_/B VGND VGND VPWR VPWR _20982_/Y sky130_fd_sc_hd__nor2_4
XFILLER_38_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22561__A1 _21105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22721_ _22796_/B VGND VGND VPWR VPWR _22722_/B sky130_fd_sc_hd__buf_2
XFILLER_53_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25440_ _25425_/CLK _25440_/D HRESETn VGND VGND VPWR VPWR _12260_/A sky130_fd_sc_hd__dfrtp_4
X_22652_ _21529_/X _22651_/X _21532_/X _24855_/Q _21533_/X VGND VGND VPWR VPWR _22653_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25433__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21603_ _21629_/A _19792_/Y VGND VGND VPWR VPWR _21605_/B sky130_fd_sc_hd__or2_4
XFILLER_16_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25371_ _25374_/CLK _25371_/D HRESETn VGND VGND VPWR VPWR _12752_/A sky130_fd_sc_hd__dfrtp_4
X_22583_ _22583_/A _16373_/A VGND VGND VPWR VPWR _22583_/X sky130_fd_sc_hd__or2_4
XANTENNA__16355__A _16355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21534_ _21529_/X _21531_/X _21532_/X _24705_/Q _21533_/X VGND VGND VPWR VPWR _21534_/X
+ sky130_fd_sc_hd__a32o_4
X_24322_ _24322_/CLK _24322_/D HRESETn VGND VGND VPWR VPWR _20990_/B sky130_fd_sc_hd__dfstp_4
XFILLER_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24253_ _24346_/CLK _17865_/Y HRESETn VGND VGND VPWR VPWR _24253_/Q sky130_fd_sc_hd__dfrtp_4
X_21465_ _21465_/A _19966_/Y VGND VGND VPWR VPWR _21467_/B sky130_fd_sc_hd__or2_4
XANTENNA__15751__B1 _24854_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22616__A2 _22534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23204_ _15090_/A _23327_/B VGND VGND VPWR VPWR _23204_/X sky130_fd_sc_hd__or2_4
X_20416_ _23371_/Q VGND VGND VPWR VPWR _20416_/Y sky130_fd_sc_hd__inv_2
X_24184_ _24373_/CLK _18375_/X HRESETn VGND VGND VPWR VPWR _24184_/Q sky130_fd_sc_hd__dfrtp_4
X_21396_ _21381_/A _20268_/Y VGND VGND VPWR VPWR _21396_/X sky130_fd_sc_hd__or2_4
XFILLER_119_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17186__A _23072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23135_ _24458_/Q _22998_/X _22885_/X VGND VGND VPWR VPWR _23135_/X sky130_fd_sc_hd__o21a_4
X_20347_ _23400_/Q VGND VGND VPWR VPWR _20347_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24386__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23066_ _23002_/A _23066_/B _23066_/C _23066_/D VGND VGND VPWR VPWR _23066_/X sky130_fd_sc_hd__or4_4
X_20278_ _20290_/A VGND VGND VPWR VPWR _20278_/X sky130_fd_sc_hd__buf_2
XFILLER_62_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24315__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22017_ _22024_/A _19935_/Y VGND VGND VPWR VPWR _22018_/C sky130_fd_sc_hd__or2_4
XFILLER_88_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13219__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_1_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23329__B1 _22797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20340__A _20339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_56_0_HCLK clkbuf_6_28_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__17008__B1 _24723_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14770_ _16173_/A _14770_/B _14555_/B VGND VGND VPWR VPWR _14781_/B sky130_fd_sc_hd__and3_4
XANTENNA__21155__B _15852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11982_ _11654_/C _11981_/X _11979_/X VGND VGND VPWR VPWR _25485_/D sky130_fd_sc_hd__o21a_4
X_23968_ _23964_/CLK _23968_/D HRESETn VGND VGND VPWR VPWR _23968_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_57_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22552__A1 _22476_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22552__B2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13721_ _13721_/A VGND VGND VPWR VPWR _13721_/X sky130_fd_sc_hd__buf_2
X_22919_ _13119_/D _21278_/X _13649_/D _21302_/X VGND VGND VPWR VPWR _22919_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23899_ _23905_/CLK _18950_/X VGND VGND VPWR VPWR _13222_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_32_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23950__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16440_ _16439_/Y _16437_/X _16359_/X _16437_/X VGND VGND VPWR VPWR _16440_/X sky130_fd_sc_hd__a2bb2o_4
X_13652_ _24030_/Q _21209_/A VGND VGND VPWR VPWR _13653_/B sky130_fd_sc_hd__nor2_4
XFILLER_44_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14242__B1 _13810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22267__A _22267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12603_ _12664_/A VGND VGND VPWR VPWR _12657_/A sky130_fd_sc_hd__buf_2
XFILLER_125_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16371_ _16371_/A _22441_/A VGND VGND VPWR VPWR _16371_/X sky130_fd_sc_hd__or2_4
XANTENNA__25103__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ _13580_/Y _14570_/A _21952_/A _13582_/Y VGND VGND VPWR VPWR _13583_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16265__A _21322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18110_ _17973_/X _18110_/B VGND VGND VPWR VPWR _18112_/B sky130_fd_sc_hd__or2_4
XFILLER_13_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15322_ _15322_/A _15322_/B VGND VGND VPWR VPWR _15322_/X sky130_fd_sc_hd__or2_4
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _25407_/Q _12533_/A _12609_/A _12533_/Y VGND VGND VPWR VPWR _12534_/X sky130_fd_sc_hd__o22a_4
X_19090_ _19090_/A VGND VGND VPWR VPWR _22060_/B sky130_fd_sc_hd__inv_2
XFILLER_125_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18041_ _18202_/A VGND VGND VPWR VPWR _18185_/A sky130_fd_sc_hd__buf_2
X_15253_ _14885_/A _15253_/B VGND VGND VPWR VPWR _15253_/X sky130_fd_sc_hd__or2_4
X_12465_ _12235_/X _12459_/X _12412_/A _12461_/Y VGND VGND VPWR VPWR _12465_/X sky130_fd_sc_hd__a211o_4
X_14204_ _20500_/A _14199_/X _13837_/X _14201_/X VGND VGND VPWR VPWR _14204_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21815__B1 _21493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12396_ _12396_/A VGND VGND VPWR VPWR _12396_/Y sky130_fd_sc_hd__inv_2
X_15184_ _15072_/B _15165_/B VGND VGND VPWR VPWR _15185_/A sky130_fd_sc_hd__or2_4
X_14135_ _14117_/C _14103_/B _14117_/C _14103_/B VGND VGND VPWR VPWR _14135_/X sky130_fd_sc_hd__a2bb2o_4
X_19992_ _19992_/A VGND VGND VPWR VPWR _19992_/X sky130_fd_sc_hd__buf_2
XFILLER_4_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14066_ _14076_/A VGND VGND VPWR VPWR _14066_/X sky130_fd_sc_hd__buf_2
X_18943_ _18942_/Y _18937_/X _17443_/X _18937_/A VGND VGND VPWR VPWR _18943_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24056__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13017_ _12306_/Y _12999_/X _13023_/A _13017_/D VGND VGND VPWR VPWR _13017_/X sky130_fd_sc_hd__or4_4
X_18874_ _18874_/A _18874_/B VGND VGND VPWR VPWR _18875_/B sky130_fd_sc_hd__or2_4
X_17825_ _17825_/A VGND VGND VPWR VPWR _17826_/B sky130_fd_sc_hd__inv_2
XANTENNA__16839__A1_N _14900_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17756_ _17756_/A _17755_/Y _16900_/Y _16941_/Y VGND VGND VPWR VPWR _17759_/C sky130_fd_sc_hd__or4_4
XANTENNA__21065__B _21017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14968_ _15249_/A _24405_/Q _25023_/Q _14967_/Y VGND VGND VPWR VPWR _14974_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21346__A2 _16453_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16707_ _16645_/A VGND VGND VPWR VPWR _16707_/X sky130_fd_sc_hd__buf_2
XFILLER_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13919_ _24957_/Q VGND VGND VPWR VPWR _13919_/X sky130_fd_sc_hd__buf_2
X_17687_ _17686_/X VGND VGND VPWR VPWR _24282_/D sky130_fd_sc_hd__inv_2
X_14899_ _15219_/C _16823_/A _15067_/D _16823_/A VGND VGND VPWR VPWR _14910_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19426_ _19017_/X VGND VGND VPWR VPWR _19426_/X sky130_fd_sc_hd__buf_2
X_16638_ _16172_/B _16624_/X VGND VGND VPWR VPWR _16638_/X sky130_fd_sc_hd__and2_4
XFILLER_63_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21081__A _23069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19357_ _19353_/Y _19356_/X _19313_/X _19356_/X VGND VGND VPWR VPWR _19357_/X sky130_fd_sc_hd__a2bb2o_4
X_16569_ _24523_/Q VGND VGND VPWR VPWR _16569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15981__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19172__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18308_ _18307_/X VGND VGND VPWR VPWR _21478_/A sky130_fd_sc_hd__buf_2
XFILLER_31_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19288_ _19287_/Y VGND VGND VPWR VPWR _19288_/X sky130_fd_sc_hd__buf_2
XANTENNA__24897__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18239_ _18235_/X _18237_/X _11803_/X _24227_/Q _18238_/X VGND VGND VPWR VPWR _24227_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_15_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15733__B1 _11778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24826__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21250_ _21250_/A _21248_/X _21250_/C VGND VGND VPWR VPWR _21250_/X sky130_fd_sc_hd__and3_4
XFILLER_102_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20201_ _21749_/B _20196_/X _19790_/A _20196_/X VGND VGND VPWR VPWR _20201_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21181_ _24199_/Q _21181_/B VGND VGND VPWR VPWR _21181_/X sky130_fd_sc_hd__or2_4
XFILLER_116_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20132_ _20132_/A VGND VGND VPWR VPWR _22071_/B sky130_fd_sc_hd__inv_2
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15238__B _15165_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20063_ _19683_/A VGND VGND VPWR VPWR _20065_/A sky130_fd_sc_hd__buf_2
X_24940_ _24643_/CLK _24940_/D HRESETn VGND VGND VPWR VPWR _24940_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24871_ _25397_/CLK _15719_/X HRESETn VGND VGND VPWR VPWR _24871_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23822_ _25044_/CLK _23822_/D VGND VGND VPWR VPWR _19169_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20965_ _12149_/X _20965_/B VGND VGND VPWR VPWR _20965_/X sky130_fd_sc_hd__and2_4
XFILLER_54_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23753_ _23772_/CLK _23753_/D VGND VGND VPWR VPWR _23753_/Q sky130_fd_sc_hd__dfxtp_4
X_22704_ _24717_/Q _22407_/B _21103_/A _22703_/X VGND VGND VPWR VPWR _22704_/X sky130_fd_sc_hd__a211o_4
X_20896_ _24047_/Q VGND VGND VPWR VPWR _20896_/Y sky130_fd_sc_hd__inv_2
X_23684_ _23683_/CLK _19563_/X VGND VGND VPWR VPWR _23684_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22087__A _23085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25423_ _25368_/CLK _12501_/X HRESETn VGND VGND VPWR VPWR _12263_/A sky130_fd_sc_hd__dfrtp_4
X_22635_ _22827_/A _22633_/X _22103_/X _22634_/X VGND VGND VPWR VPWR _22636_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22837__A2 _22833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15972__B1 _24748_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19163__B1 _19071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25354_ _25354_/CLK _25354_/D HRESETn VGND VGND VPWR VPWR _21006_/A sky130_fd_sc_hd__dfrtp_4
X_22566_ _16898_/X _22425_/A _12282_/C _22489_/A VGND VGND VPWR VPWR _22566_/X sky130_fd_sc_hd__o22a_4
X_21517_ _23100_/A VGND VGND VPWR VPWR _23306_/A sky130_fd_sc_hd__buf_2
XANTENNA__16623__A2_N _16545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24305_ _24305_/CLK _24305_/D HRESETn VGND VGND VPWR VPWR _17605_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_6_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15724__B1 _24868_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22497_ _22441_/X _22494_/X _22444_/X _22496_/X VGND VGND VPWR VPWR _22498_/B sky130_fd_sc_hd__o22a_4
X_25285_ _25478_/CLK _13674_/X HRESETn VGND VGND VPWR VPWR _25285_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24567__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12250_ _12249_/X _24750_/Q _12249_/X _24750_/Q VGND VGND VPWR VPWR _12250_/X sky130_fd_sc_hd__a2bb2o_4
X_21448_ _21455_/A VGND VGND VPWR VPWR _21449_/A sky130_fd_sc_hd__buf_2
X_24236_ _23826_/CLK _24236_/D HRESETn VGND VGND VPWR VPWR _24236_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20335__A _20335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12181_ _22267_/A VGND VGND VPWR VPWR _12181_/Y sky130_fd_sc_hd__inv_2
X_24167_ _24502_/CLK _18520_/Y HRESETn VGND VGND VPWR VPWR _24167_/Q sky130_fd_sc_hd__dfrtp_4
X_21379_ _21377_/A VGND VGND VPWR VPWR _21398_/A sky130_fd_sc_hd__buf_2
XFILLER_135_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23118_ _22782_/A VGND VGND VPWR VPWR _23124_/A sky130_fd_sc_hd__buf_2
XANTENNA__23014__A2 _21287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24098_ _23933_/CLK _20963_/X HRESETn VGND VGND VPWR VPWR _12127_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_27_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22550__A _22550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15940_ HWDATA[29] VGND VGND VPWR VPWR _15940_/X sky130_fd_sc_hd__buf_2
XANTENNA__19565__A2_N _19562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23049_ _17257_/A _22908_/X _12896_/A _22909_/X VGND VGND VPWR VPWR _23049_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21576__A2 _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15871_ _12820_/Y _15869_/X _11754_/X _15869_/X VGND VGND VPWR VPWR _15871_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12788__A _24774_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17610_ _17609_/X VGND VGND VPWR VPWR _17610_/Y sky130_fd_sc_hd__inv_2
X_14822_ _14870_/B VGND VGND VPWR VPWR _14880_/B sky130_fd_sc_hd__buf_2
XANTENNA__15164__A _15171_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18590_ _18418_/Y _18585_/X VGND VGND VPWR VPWR _18591_/B sky130_fd_sc_hd__nand2_4
XANTENNA__25355__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21328__A2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17541_ _24298_/Q VGND VGND VPWR VPWR _17541_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14753_ _14750_/X VGND VGND VPWR VPWR _14753_/Y sky130_fd_sc_hd__inv_2
X_11965_ _11964_/X VGND VGND VPWR VPWR _11965_/X sky130_fd_sc_hd__buf_2
XFILLER_17_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13704_ _13699_/X _13680_/X _13702_/Y _13703_/X _13693_/C VGND VGND VPWR VPWR _13704_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_45_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_143_0_HCLK clkbuf_7_71_0_HCLK/X VGND VGND VPWR VPWR _24197_/CLK sky130_fd_sc_hd__clkbuf_1
X_17472_ _17472_/A _17472_/B VGND VGND VPWR VPWR _17472_/Y sky130_fd_sc_hd__nor2_4
XFILLER_72_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14684_ _14684_/A VGND VGND VPWR VPWR _14746_/A sky130_fd_sc_hd__inv_2
XANTENNA__14215__B1 _13810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11896_ _11900_/A VGND VGND VPWR VPWR _11896_/X sky130_fd_sc_hd__buf_2
XANTENNA__15558__A3 _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15412__C1 _15339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19211_ _19197_/X VGND VGND VPWR VPWR _19211_/X sky130_fd_sc_hd__buf_2
X_16423_ _22608_/A VGND VGND VPWR VPWR _16423_/Y sky130_fd_sc_hd__inv_2
X_13635_ _13635_/A _13598_/X VGND VGND VPWR VPWR _13635_/X sky130_fd_sc_hd__or2_4
XFILLER_73_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19503__A2_N _19500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15963__B1 _15962_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22828__A2 _22790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19142_ _19141_/Y _19137_/X _19117_/X _19137_/X VGND VGND VPWR VPWR _19142_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16354_ _21852_/A VGND VGND VPWR VPWR _16354_/Y sky130_fd_sc_hd__inv_2
X_13566_ _13566_/A VGND VGND VPWR VPWR _14561_/A sky130_fd_sc_hd__inv_2
XFILLER_125_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22725__A _22574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24990__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15305_ _15133_/Y _15128_/Y _15305_/C VGND VGND VPWR VPWR _15336_/B sky130_fd_sc_hd__or3_4
X_12517_ _25413_/Q VGND VGND VPWR VPWR _12517_/Y sky130_fd_sc_hd__inv_2
X_19073_ _13337_/B VGND VGND VPWR VPWR _19073_/Y sky130_fd_sc_hd__inv_2
X_16285_ HWDATA[30] VGND VGND VPWR VPWR _16285_/X sky130_fd_sc_hd__buf_2
XANTENNA__15715__B1 _24872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13497_ _13497_/A VGND VGND VPWR VPWR _13497_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16723__A _16723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18024_ _18024_/A _18024_/B VGND VGND VPWR VPWR _18027_/B sky130_fd_sc_hd__or2_4
X_15236_ _15210_/B _15210_/C _15199_/X _15233_/B VGND VGND VPWR VPWR _15236_/X sky130_fd_sc_hd__a211o_4
X_12448_ _25437_/Q _12448_/B VGND VGND VPWR VPWR _12449_/C sky130_fd_sc_hd__or2_4
XANTENNA__23253__A2 _22824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20245__A _20232_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24237__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15730__A3 _15729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_11_0_HCLK_A clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11867__A _11867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15167_ _15169_/B VGND VGND VPWR VPWR _15167_/Y sky130_fd_sc_hd__inv_2
X_12379_ _12377_/Y _12296_/A _12993_/A _24810_/Q VGND VGND VPWR VPWR _12379_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14118_ _14117_/X VGND VGND VPWR VPWR _14118_/Y sky130_fd_sc_hd__inv_2
X_15098_ _24971_/Q VGND VGND VPWR VPWR _15299_/B sky130_fd_sc_hd__inv_2
X_19975_ _11922_/A VGND VGND VPWR VPWR _19975_/X sky130_fd_sc_hd__buf_2
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17554__A _17837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14049_ _14006_/A _14047_/Y _14001_/D _14049_/D VGND VGND VPWR VPWR _14049_/X sky130_fd_sc_hd__and4_4
X_18926_ _18921_/Y _18925_/X _17418_/X _18925_/X VGND VGND VPWR VPWR _23908_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23275__B _21519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18968__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18857_ _16503_/Y _18688_/A _16503_/Y _18688_/A VGND VGND VPWR VPWR _18857_/X sky130_fd_sc_hd__a2bb2o_4
X_17808_ _17759_/A _17753_/Y _17792_/C _17751_/X VGND VGND VPWR VPWR _17830_/B sky130_fd_sc_hd__or4_4
XANTENNA__23308__A3 _21514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18788_ _18788_/A VGND VGND VPWR VPWR _18788_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25096__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13257__B2 _11965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21319__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17739_ _24275_/Q VGND VGND VPWR VPWR _17765_/C sky130_fd_sc_hd__inv_2
XFILLER_36_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25025__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19393__B1 _19370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20750_ _13119_/C _20772_/C VGND VGND VPWR VPWR _20750_/X sky130_fd_sc_hd__or2_4
XFILLER_51_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14206__B1 _13840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19409_ _19406_/Y _19401_/X _19407_/X _19408_/X VGND VGND VPWR VPWR _23738_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20681_ _15638_/Y _20677_/X _23997_/Q _20680_/X VGND VGND VPWR VPWR _20681_/X sky130_fd_sc_hd__o22a_4
XFILLER_56_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14418__A _16528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19145__B1 _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22420_ _22419_/X VGND VGND VPWR VPWR _22424_/A sky130_fd_sc_hd__buf_2
XFILLER_31_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22351_ _17722_/A _22350_/X _17728_/A VGND VGND VPWR VPWR _22351_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24660__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21302_ _21302_/A VGND VGND VPWR VPWR _21302_/X sky130_fd_sc_hd__buf_2
X_25070_ _25070_/CLK _25070_/D HRESETn VGND VGND VPWR VPWR _25070_/Q sky130_fd_sc_hd__dfrtp_4
X_22282_ _22278_/X _22279_/X _22280_/X _22281_/X VGND VGND VPWR VPWR _22283_/B sky130_fd_sc_hd__o22a_4
XANTENNA__23244__A2 _22393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17448__B _17447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13193__B1 _11958_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24021_ _24049_/CLK _20785_/X HRESETn VGND VGND VPWR VPWR _24021_/Q sky130_fd_sc_hd__dfrtp_4
X_21233_ _14710_/Y VGND VGND VPWR VPWR _21233_/X sky130_fd_sc_hd__buf_2
XFILLER_102_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11777__A _11777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21164_ _21173_/A _21164_/B VGND VGND VPWR VPWR _21164_/X sky130_fd_sc_hd__or2_4
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22370__A _21616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20115_ _20115_/A VGND VGND VPWR VPWR _21756_/B sky130_fd_sc_hd__inv_2
X_21095_ _21306_/A VGND VGND VPWR VPWR _21095_/X sky130_fd_sc_hd__buf_2
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22755__A1 _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20046_ _22368_/B _20045_/X _19777_/X _20045_/X VGND VGND VPWR VPWR _20046_/X sky130_fd_sc_hd__a2bb2o_4
X_24923_ _24923_/CLK _15520_/X HRESETn VGND VGND VPWR VPWR _11730_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24854_ _24865_/CLK _15751_/X HRESETn VGND VGND VPWR VPWR _24854_/Q sky130_fd_sc_hd__dfrtp_4
X_23805_ _23805_/CLK _19217_/X VGND VGND VPWR VPWR _18222_/B sky130_fd_sc_hd__dfxtp_4
X_24785_ _24785_/CLK _24785_/D HRESETn VGND VGND VPWR VPWR _22651_/A sky130_fd_sc_hd__dfrtp_4
X_21997_ _21978_/C _22389_/B VGND VGND VPWR VPWR _21997_/Y sky130_fd_sc_hd__nor2_4
XPHY_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18726__C _18743_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11750_/A VGND VGND VPWR VPWR _11777_/A sky130_fd_sc_hd__buf_2
XANTENNA__16198__B1 _15944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21433__B _22590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23736_ _23718_/CLK _19413_/X VGND VGND VPWR VPWR _19412_/A sky130_fd_sc_hd__dfxtp_4
X_20948_ _20946_/Y _20947_/Y _13667_/X VGND VGND VPWR VPWR _20948_/X sky130_fd_sc_hd__o21a_4
XFILLER_121_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_216_0_HCLK clkbuf_8_217_0_HCLK/A VGND VGND VPWR VPWR _24055_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _25278_/Q _24223_/Q _13690_/A _22532_/A VGND VGND VPWR VPWR _11688_/B sky130_fd_sc_hd__o22a_4
XPHY_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23667_ _23623_/CLK _23667_/D VGND VGND VPWR VPWR _23667_/Q sky130_fd_sc_hd__dfxtp_4
X_20879_ _20879_/A _20879_/B VGND VGND VPWR VPWR _20879_/X sky130_fd_sc_hd__or2_4
XANTENNA__24748__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12261__A2_N _12259_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13452_/A _23654_/Q VGND VGND VPWR VPWR _13421_/C sky130_fd_sc_hd__or2_4
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25406_ _25400_/CLK _25406_/D HRESETn VGND VGND VPWR VPWR _25406_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22618_ _22617_/X VGND VGND VPWR VPWR _22618_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22286__A3 _22396_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23598_ _23598_/CLK _23598_/D VGND VGND VPWR VPWR _19817_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17698__B1 _17601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13351_ _13297_/X _13343_/X _13351_/C VGND VGND VPWR VPWR _13351_/X sky130_fd_sc_hd__and3_4
XFILLER_128_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25337_ _24852_/CLK _13067_/X HRESETn VGND VGND VPWR VPWR _25337_/Q sky130_fd_sc_hd__dfrtp_4
X_22549_ _22549_/A _22549_/B VGND VGND VPWR VPWR _22549_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__16543__A _16795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12302_ _12302_/A VGND VGND VPWR VPWR _12303_/A sky130_fd_sc_hd__inv_2
XFILLER_127_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16070_ _16069_/Y _16067_/X _15474_/X _16067_/X VGND VGND VPWR VPWR _16070_/X sky130_fd_sc_hd__a2bb2o_4
X_13282_ _13387_/A _13282_/B VGND VGND VPWR VPWR _13282_/X sky130_fd_sc_hd__or2_4
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25268_ _24252_/CLK _13733_/X HRESETn VGND VGND VPWR VPWR _25268_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24330__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15712__A3 _15553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15021_ _15014_/X _15016_/X _15021_/C _15021_/D VGND VGND VPWR VPWR _15021_/X sky130_fd_sc_hd__or4_4
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17493__A1_N _11706_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12233_ _12280_/A _12231_/Y _25425_/Q _12232_/Y VGND VGND VPWR VPWR _12240_/B sky130_fd_sc_hd__a2bb2o_4
X_24219_ _24219_/CLK _24219_/D HRESETn VGND VGND VPWR VPWR _24219_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25199_ _25199_/CLK _25199_/D HRESETn VGND VGND VPWR VPWR _14098_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22994__A1 _24523_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12164_ _18370_/A _12159_/X _12163_/X VGND VGND VPWR VPWR _25455_/D sky130_fd_sc_hd__a21o_4
XFILLER_107_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22280__A _22280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12095_ _12095_/A VGND VGND VPWR VPWR _12095_/Y sky130_fd_sc_hd__inv_2
X_16972_ _24379_/Q VGND VGND VPWR VPWR _16972_/Y sky130_fd_sc_hd__inv_2
X_19760_ _19757_/Y _19752_/X _19758_/X _19759_/X VGND VGND VPWR VPWR _23618_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25536__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22746__B2 _22922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15923_ _15843_/A _15925_/B VGND VGND VPWR VPWR _15923_/X sky130_fd_sc_hd__or2_4
X_18711_ _18711_/A VGND VGND VPWR VPWR _18712_/B sky130_fd_sc_hd__inv_2
XFILLER_7_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19691_ _19689_/Y _19685_/X _19645_/X _19690_/X VGND VGND VPWR VPWR _19691_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18642_ _16620_/A _18639_/Y _16611_/A _18786_/C VGND VGND VPWR VPWR _18642_/X sky130_fd_sc_hd__a2bb2o_4
X_15854_ _22835_/A VGND VGND VPWR VPWR _15854_/X sky130_fd_sc_hd__buf_2
XFILLER_91_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_26_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_14805_ _14805_/A VGND VGND VPWR VPWR _14820_/A sky130_fd_sc_hd__inv_2
X_18573_ _18469_/B _18576_/B VGND VGND VPWR VPWR _18573_/Y sky130_fd_sc_hd__nand2_4
X_15785_ _15931_/A VGND VGND VPWR VPWR _15925_/B sky130_fd_sc_hd__buf_2
XFILLER_91_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12997_ _12352_/Y _12347_/Y _13071_/B VGND VGND VPWR VPWR _13043_/B sky130_fd_sc_hd__or3_4
XANTENNA__19375__B1 _19307_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17524_ _17497_/X _17505_/X _17514_/X _17523_/X VGND VGND VPWR VPWR _17524_/X sky130_fd_sc_hd__or4_4
X_14736_ _14736_/A VGND VGND VPWR VPWR _14736_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11948_ _11948_/A VGND VGND VPWR VPWR _11948_/X sky130_fd_sc_hd__buf_2
XFILLER_73_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17455_ _24197_/Q _13177_/A _20231_/C _13177_/Y VGND VGND VPWR VPWR _17457_/A sky130_fd_sc_hd__o22a_4
X_14667_ _13624_/A _19038_/C _14659_/B VGND VGND VPWR VPWR _14667_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15936__B1 _24765_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11879_ _11700_/X _11879_/B VGND VGND VPWR VPWR _11899_/A sky130_fd_sc_hd__or2_4
XANTENNA__24489__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16406_ _16389_/A VGND VGND VPWR VPWR _16406_/X sky130_fd_sc_hd__buf_2
X_13618_ _25058_/Q VGND VGND VPWR VPWR _13618_/Y sky130_fd_sc_hd__inv_2
X_17386_ _23982_/Q VGND VGND VPWR VPWR _17387_/A sky130_fd_sc_hd__inv_2
XFILLER_60_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14598_ _14598_/A _14564_/X VGND VGND VPWR VPWR _14598_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24418__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22455__A _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15951__A3 HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19125_ _19124_/Y _19120_/X _19010_/X _19106_/Y VGND VGND VPWR VPWR _19125_/X sky130_fd_sc_hd__a2bb2o_4
X_16337_ _16324_/A VGND VGND VPWR VPWR _16337_/X sky130_fd_sc_hd__buf_2
X_13549_ _21952_/A VGND VGND VPWR VPWR _13549_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11973__A1 _21504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19056_ _19055_/X VGND VGND VPWR VPWR _19056_/X sky130_fd_sc_hd__buf_2
XANTENNA__11973__B2 _13678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16268_ _16268_/A VGND VGND VPWR VPWR _16268_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24071__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18007_ _18087_/A VGND VGND VPWR VPWR _18184_/A sky130_fd_sc_hd__buf_2
X_15219_ _15219_/A _15219_/B _15219_/C _15211_/B VGND VGND VPWR VPWR _15219_/X sky130_fd_sc_hd__or4_4
X_16199_ _23165_/A VGND VGND VPWR VPWR _16199_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24000__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12922__B1 _12874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19958_ _22016_/B _19952_/X _19618_/X _19957_/X VGND VGND VPWR VPWR _23546_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25277__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_108_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_217_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18909_ _18909_/A VGND VGND VPWR VPWR _18909_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25206__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19889_ _19889_/A VGND VGND VPWR VPWR _19902_/A sky130_fd_sc_hd__inv_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21920_ _21942_/A _21920_/B VGND VGND VPWR VPWR _21921_/C sky130_fd_sc_hd__or2_4
XFILLER_95_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21851_ _21019_/A VGND VGND VPWR VPWR _22406_/B sky130_fd_sc_hd__buf_2
XANTENNA__20917__A1_N _20909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20802_ _20680_/X _20801_/Y _24908_/Q _20725_/X VGND VGND VPWR VPWR _24025_/D sky130_fd_sc_hd__a2bb2o_4
X_21782_ _21816_/B _21780_/X _21502_/A _21781_/X VGND VGND VPWR VPWR _21782_/X sky130_fd_sc_hd__a211o_4
XFILLER_23_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24570_ _24465_/CLK _16440_/X HRESETn VGND VGND VPWR VPWR _24570_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23521_ _24923_/CLK _23521_/D VGND VGND VPWR VPWR _23521_/Q sky130_fd_sc_hd__dfxtp_4
X_20733_ _20721_/X _20732_/Y _24892_/Q _20726_/X VGND VGND VPWR VPWR _20733_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20920__B1 _20845_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19118__B1 _19117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24841__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20664_ _20664_/A _20474_/B VGND VGND VPWR VPWR _20665_/C sky130_fd_sc_hd__or2_4
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23452_ _23446_/CLK _23452_/D VGND VGND VPWR VPWR _20209_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_46_0_HCLK clkbuf_8_47_0_HCLK/A VGND VGND VPWR VPWR _25488_/CLK sky130_fd_sc_hd__clkbuf_1
X_22403_ _22271_/X _22402_/X _21290_/C _24710_/Q _21067_/X VGND VGND VPWR VPWR _22403_/X
+ sky130_fd_sc_hd__a32o_4
X_23383_ _24219_/CLK _23383_/D VGND VGND VPWR VPWR _23383_/Q sky130_fd_sc_hd__dfxtp_4
X_20595_ _20428_/B VGND VGND VPWR VPWR _20595_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22084__B _23082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25122_ _25122_/CLK _25122_/D HRESETn VGND VGND VPWR VPWR _25122_/Q sky130_fd_sc_hd__dfstp_4
X_22334_ _21917_/X _22332_/X _22333_/X VGND VGND VPWR VPWR _22334_/X sky130_fd_sc_hd__and3_4
XFILLER_87_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22265_ _21570_/X VGND VGND VPWR VPWR _22265_/X sky130_fd_sc_hd__buf_2
X_25053_ _25054_/CLK _25053_/D HRESETn VGND VGND VPWR VPWR _22036_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_30_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22812__B _22810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21216_ _15665_/A _21215_/X _13671_/Y _15665_/A VGND VGND VPWR VPWR _21216_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12913__B1 _12866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24004_ _24035_/CLK _24004_/D HRESETn VGND VGND VPWR VPWR _13129_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16104__B1 _11764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22196_ _14712_/A _22191_/X _22195_/X VGND VGND VPWR VPWR _22196_/X sky130_fd_sc_hd__or3_4
X_21147_ _21350_/B _21146_/X _21116_/A VGND VGND VPWR VPWR _21147_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15707__A _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17194__A _23246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21078_ _15852_/Y VGND VGND VPWR VPWR _21859_/C sky130_fd_sc_hd__buf_2
XFILLER_101_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12920_ _12810_/A _12919_/Y VGND VGND VPWR VPWR _12920_/X sky130_fd_sc_hd__or2_4
X_20029_ _20036_/A VGND VGND VPWR VPWR _20029_/X sky130_fd_sc_hd__buf_2
XANTENNA__13227__A _13227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24906_ _24055_/CLK _15573_/X HRESETn VGND VGND VPWR VPWR _15572_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14948__A2_N _24413_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12851_ _12806_/A _12799_/A _12849_/X _12851_/D VGND VGND VPWR VPWR _12852_/B sky130_fd_sc_hd__or4_4
XFILLER_73_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24837_ _24830_/CLK _24837_/D HRESETn VGND VGND VPWR VPWR _24837_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11970__A _11958_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19357__B1 _19313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24929__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11802_ _11802_/A VGND VGND VPWR VPWR _11802_/Y sky130_fd_sc_hd__inv_2
X_15570_ _15570_/A VGND VGND VPWR VPWR _15570_/Y sky130_fd_sc_hd__inv_2
X_12782_ _24801_/Q VGND VGND VPWR VPWR _12782_/Y sky130_fd_sc_hd__inv_2
XPHY_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24768_ _24806_/CLK _15926_/X HRESETn VGND VGND VPWR VPWR _12983_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _23951_/Q VGND VGND VPWR VPWR _14521_/X sky130_fd_sc_hd__buf_2
XANTENNA__22900__B2 _22480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11733_ _11733_/A _21027_/A VGND VGND VPWR VPWR _11734_/A sky130_fd_sc_hd__or2_4
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23719_ _23887_/CLK _19460_/X VGND VGND VPWR VPWR _19458_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_15_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24582__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24699_ _24699_/CLK _16089_/X HRESETn VGND VGND VPWR VPWR _23310_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22438__A1_N _17350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17240_ _17240_/A VGND VGND VPWR VPWR _17240_/Y sky130_fd_sc_hd__inv_2
XPHY_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14381_/A VGND VGND VPWR VPWR _14452_/X sky130_fd_sc_hd__buf_2
XPHY_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11664_/A VGND VGND VPWR VPWR _11664_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16591__B1 _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24511__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _13260_/X _13403_/B _13403_/C VGND VGND VPWR VPWR _13403_/X sky130_fd_sc_hd__and3_4
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17171_ _16299_/Y _17295_/A _16299_/Y _17295_/A VGND VGND VPWR VPWR _17171_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14383_ _14383_/A VGND VGND VPWR VPWR _14384_/A sky130_fd_sc_hd__buf_2
XFILLER_10_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16122_ _16122_/A VGND VGND VPWR VPWR _16122_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20507__B _14207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _13200_/X _13315_/X _13333_/X _25318_/Q _11965_/X VGND VGND VPWR VPWR _13334_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_122_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16053_ _16051_/Y _16047_/X _15756_/X _16052_/X VGND VGND VPWR VPWR _16053_/X sky130_fd_sc_hd__a2bb2o_4
X_13265_ _13379_/A _13265_/B VGND VGND VPWR VPWR _13265_/X sky130_fd_sc_hd__or2_4
X_15004_ _25011_/Q _15003_/A _15219_/C _15003_/Y VGND VGND VPWR VPWR _15004_/X sky130_fd_sc_hd__o22a_4
X_12216_ _12399_/A VGND VGND VPWR VPWR _12385_/A sky130_fd_sc_hd__inv_2
X_13196_ _13195_/X VGND VGND VPWR VPWR _13196_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22431__A3 _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19812_ _13363_/B VGND VGND VPWR VPWR _19812_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17843__B1 _17790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_HCLK_A HCLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12147_ _24100_/Q _12147_/B VGND VGND VPWR VPWR _12148_/A sky130_fd_sc_hd__and2_4
XFILLER_97_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15617__A _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25370__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19743_ _19729_/Y VGND VGND VPWR VPWR _19743_/X sky130_fd_sc_hd__buf_2
XANTENNA__15336__B _15336_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12078_ _25471_/Q VGND VGND VPWR VPWR _12078_/Y sky130_fd_sc_hd__inv_2
X_16955_ _17805_/A VGND VGND VPWR VPWR _16955_/X sky130_fd_sc_hd__buf_2
XANTENNA__19596__B1 _19547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17254__D _17253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15906_ _15705_/X _15894_/X _15836_/X _24776_/Q _15864_/A VGND VGND VPWR VPWR _15906_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16886_ _16884_/Y _16880_/X _16885_/X _16880_/X VGND VGND VPWR VPWR _16886_/X sky130_fd_sc_hd__a2bb2o_4
X_19674_ _19673_/Y _19669_/X _19599_/X _19669_/X VGND VGND VPWR VPWR _19674_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15837_ _15824_/X _15835_/X _15836_/X _24811_/Q _15793_/A VGND VGND VPWR VPWR _15837_/X
+ sky130_fd_sc_hd__a32o_4
X_18625_ _18625_/A _18620_/X _18625_/C _18624_/X VGND VGND VPWR VPWR _18636_/C sky130_fd_sc_hd__or4_4
XANTENNA__12976__A _12976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16448__A _16448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11880__A _11700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21073__B _21073_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15768_ _18254_/A VGND VGND VPWR VPWR _15768_/X sky130_fd_sc_hd__buf_2
X_18556_ _18468_/Y _18550_/X _18552_/Y _18487_/X VGND VGND VPWR VPWR _18556_/X sky130_fd_sc_hd__a211o_4
XFILLER_45_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14719_ _14719_/A _14719_/B _14713_/X _14718_/X VGND VGND VPWR VPWR _14719_/X sky130_fd_sc_hd__or4_4
X_17507_ _25526_/Q _24297_/Q _11783_/Y _17567_/A VGND VGND VPWR VPWR _17514_/A sky130_fd_sc_hd__o22a_4
X_18487_ _18821_/B VGND VGND VPWR VPWR _18487_/X sky130_fd_sc_hd__buf_2
XANTENNA__15909__B1 _15840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15699_ _15681_/A _15698_/X _15690_/X VGND VGND VPWR VPWR _15699_/X sky130_fd_sc_hd__o21a_4
X_17438_ _24312_/Q VGND VGND VPWR VPWR _17438_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24252__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_5_0_HCLK clkbuf_8_5_0_HCLK/A VGND VGND VPWR VPWR _23846_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_53_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17369_ _17369_/A _17369_/B VGND VGND VPWR VPWR _17369_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__16183__A _16183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19108_ _19104_/Y _19107_/X _19018_/X _19107_/X VGND VGND VPWR VPWR _23844_/D sky130_fd_sc_hd__a2bb2o_4
X_20380_ _18230_/B _19535_/X VGND VGND VPWR VPWR _20380_/X sky130_fd_sc_hd__or2_4
XANTENNA__22913__A _22913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19039_ _19038_/X VGND VGND VPWR VPWR _19052_/A sky130_fd_sc_hd__buf_2
XANTENNA__12216__A _12399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25458__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22050_ _21245_/A VGND VGND VPWR VPWR _22050_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21529__A _21108_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21001_ sda_oen_o_S5 _24937_/Q _20996_/A _15426_/X _21000_/Y VGND VGND VPWR VPWR
+ _21001_/X sky130_fd_sc_hd__a32o_4
XFILLER_138_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25040__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22952_ _23021_/A _22952_/B _22952_/C VGND VGND VPWR VPWR _22952_/X sky130_fd_sc_hd__and3_4
XFILLER_83_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15048__A2_N _24444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21903_ _14689_/A _21903_/B VGND VGND VPWR VPWR _21903_/X sky130_fd_sc_hd__or2_4
XFILLER_3_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12886__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22883_ _23170_/A VGND VGND VPWR VPWR _23065_/A sky130_fd_sc_hd__buf_2
XFILLER_102_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24622_ _24712_/CLK _24622_/D HRESETn VGND VGND VPWR VPWR _23039_/A sky130_fd_sc_hd__dfrtp_4
X_21834_ _21106_/X _21828_/Y _21547_/A _21833_/X VGND VGND VPWR VPWR _21834_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22867__A2_N _22862_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24553_ _24553_/CLK _16492_/X HRESETn VGND VGND VPWR VPWR _16490_/A sky130_fd_sc_hd__dfrtp_4
X_21765_ _21623_/A _21765_/B VGND VGND VPWR VPWR _21766_/C sky130_fd_sc_hd__or2_4
XFILLER_102_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23504_ _24208_/CLK _23504_/D VGND VGND VPWR VPWR _13348_/B sky130_fd_sc_hd__dfxtp_4
X_20716_ _20715_/X VGND VGND VPWR VPWR _20716_/Y sky130_fd_sc_hd__inv_2
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16573__B1 _16403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24484_ _24413_/CLK _24484_/D HRESETn VGND VGND VPWR VPWR _24484_/Q sky130_fd_sc_hd__dfrtp_4
X_21696_ _23306_/A _21696_/B VGND VGND VPWR VPWR _21696_/X sky130_fd_sc_hd__and2_4
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23435_ _23434_/CLK _20257_/X VGND VGND VPWR VPWR _23435_/Q sky130_fd_sc_hd__dfxtp_4
X_20647_ _20650_/B _20646_/Y _20651_/C VGND VGND VPWR VPWR _20647_/X sky130_fd_sc_hd__and3_4
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22110__A2 _22106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20578_ _18879_/A _18878_/X VGND VGND VPWR VPWR _20579_/B sky130_fd_sc_hd__nand2_4
X_23366_ _25098_/CLK scl_oen_o_S4 VGND VGND VPWR VPWR _20969_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23975__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25105_ _25113_/CLK _14484_/X HRESETn VGND VGND VPWR VPWR _14483_/A sky130_fd_sc_hd__dfrtp_4
X_22317_ _14185_/Y _14192_/X _14254_/Y _14257_/A VGND VGND VPWR VPWR _22318_/A sky130_fd_sc_hd__o22a_4
XANTENNA__25199__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23297_ _16799_/A _22135_/X _22797_/X _23296_/X VGND VGND VPWR VPWR _23298_/C sky130_fd_sc_hd__a211o_4
XFILLER_124_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13050_ _12990_/B _13045_/B _13010_/A _13047_/B VGND VGND VPWR VPWR _13050_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21439__A _11720_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25036_ _25029_/CLK _14851_/X HRESETn VGND VGND VPWR VPWR _14815_/C sky130_fd_sc_hd__dfrtp_4
X_22248_ _17720_/X _22244_/X _22248_/C VGND VGND VPWR VPWR _22248_/X sky130_fd_sc_hd__or3_4
XANTENNA__17636__B _17525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12001_ _12001_/A VGND VGND VPWR VPWR _12001_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15437__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11965__A _11964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22179_ _21332_/Y _22165_/X _22167_/X _22171_/Y _22178_/X VGND VGND VPWR VPWR _22179_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_26_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16740_ _15051_/Y _16739_/X _15723_/X _16739_/X VGND VGND VPWR VPWR _24459_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17652__A _17624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13952_ _13952_/A _13941_/Y _24954_/Q _13952_/D VGND VGND VPWR VPWR _13952_/X sky130_fd_sc_hd__and4_4
XANTENNA__14887__A2_N _24412_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12903_ _12927_/A _12924_/A _12902_/X VGND VGND VPWR VPWR _12903_/X sky130_fd_sc_hd__or3_4
X_16671_ _16664_/A VGND VGND VPWR VPWR _16671_/X sky130_fd_sc_hd__buf_2
XANTENNA__18250__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13883_ _23989_/Q _13882_/X _25172_/Q _13856_/Y VGND VGND VPWR VPWR _25231_/D sky130_fd_sc_hd__o22a_4
XFILLER_98_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12796__A _24777_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24763__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15622_ _24886_/Q VGND VGND VPWR VPWR _22281_/A sky130_fd_sc_hd__inv_2
X_18410_ _23068_/A _18409_/A _16204_/Y _18460_/B VGND VGND VPWR VPWR _18413_/C sky130_fd_sc_hd__o22a_4
XFILLER_61_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12834_ _12833_/Y _24778_/Q _12845_/A _24775_/Q VGND VGND VPWR VPWR _12835_/D sky130_fd_sc_hd__a2bb2o_4
X_19390_ _19388_/Y _19384_/X _19389_/X _19384_/X VGND VGND VPWR VPWR _19390_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18341_ _13143_/X _18340_/X _13143_/X _18340_/X VGND VGND VPWR VPWR _18341_/X sky130_fd_sc_hd__a2bb2o_4
X_15553_ HWDATA[31] VGND VGND VPWR VPWR _15553_/X sky130_fd_sc_hd__buf_2
X_12765_ _22857_/A VGND VGND VPWR VPWR _12765_/Y sky130_fd_sc_hd__inv_2
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _20441_/C _14503_/B _14502_/X _14503_/Y VGND VGND VPWR VPWR _25099_/D sky130_fd_sc_hd__a211o_4
XFILLER_128_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12814__A1_N _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11716_/A VGND VGND VPWR VPWR _15991_/C sky130_fd_sc_hd__buf_2
X_18272_ _18272_/A _18230_/B VGND VGND VPWR VPWR _18272_/X sky130_fd_sc_hd__or2_4
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15484_/A _15484_/B VGND VGND VPWR VPWR _24063_/D sky130_fd_sc_hd__nor2_4
XANTENNA__16564__B1 _16393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12570_/A _12695_/Y VGND VGND VPWR VPWR _12696_/X sky130_fd_sc_hd__or2_4
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15906__A3 _15836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17223_ _23009_/A _17222_/Y _16313_/Y _22939_/A VGND VGND VPWR VPWR _17223_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ _22316_/B VGND VGND VPWR VPWR _15462_/A sky130_fd_sc_hd__buf_2
XANTENNA__22637__B1 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _25539_/Q VGND VGND VPWR VPWR _11647_/X sky130_fd_sc_hd__buf_2
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18305__A1 _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17154_ _16993_/Y _17161_/A VGND VGND VPWR VPWR _17159_/B sky130_fd_sc_hd__or2_4
X_14366_ _25144_/Q _14348_/Y _25143_/Q _14344_/X VGND VGND VPWR VPWR _14366_/X sky130_fd_sc_hd__o22a_4
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_92_0_HCLK clkbuf_8_93_0_HCLK/A VGND VGND VPWR VPWR _24117_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_7_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22652__A3 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16105_ _16105_/A VGND VGND VPWR VPWR _16105_/Y sky130_fd_sc_hd__inv_2
X_13317_ _13317_/A _13317_/B VGND VGND VPWR VPWR _13318_/C sky130_fd_sc_hd__or2_4
XFILLER_116_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17085_ _17085_/A _17088_/B VGND VGND VPWR VPWR _17086_/C sky130_fd_sc_hd__or2_4
XFILLER_13_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21860__A1 _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14297_ _14291_/A _14301_/B _13640_/X VGND VGND VPWR VPWR _14297_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_115_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16036_ _16033_/Y _16035_/X _11796_/X _16035_/X VGND VGND VPWR VPWR _16036_/X sky130_fd_sc_hd__a2bb2o_4
X_13248_ _13248_/A VGND VGND VPWR VPWR _13452_/A sky130_fd_sc_hd__buf_2
XFILLER_83_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12353__B2 _24820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13179_ _13251_/A _23860_/Q VGND VGND VPWR VPWR _13179_/X sky130_fd_sc_hd__or2_4
XFILLER_124_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17987_ _17995_/A VGND VGND VPWR VPWR _18181_/A sky130_fd_sc_hd__buf_2
XFILLER_96_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19726_ _19725_/Y _19720_/X _19658_/X _19706_/Y VGND VGND VPWR VPWR _23629_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16938_ _16110_/Y _24267_/Q _22556_/A _16898_/X VGND VGND VPWR VPWR _16938_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21084__A _21071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19657_ _19657_/A VGND VGND VPWR VPWR _19657_/Y sky130_fd_sc_hd__inv_2
X_16869_ _16866_/Y _16859_/X _16867_/X _16868_/X VGND VGND VPWR VPWR _16869_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18608_ _18607_/Y VGND VGND VPWR VPWR _18608_/X sky130_fd_sc_hd__buf_2
XFILLER_80_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19588_ _19587_/X VGND VGND VPWR VPWR _19588_/X sky130_fd_sc_hd__buf_2
XFILLER_129_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22908__A _22419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24433__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18539_ _18541_/A _18539_/B _18538_/Y VGND VGND VPWR VPWR _18539_/X sky130_fd_sc_hd__and3_4
XANTENNA__19741__B1 _19740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21550_ _25233_/Q VGND VGND VPWR VPWR _21550_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21531__B _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20501_ _20505_/C _20500_/X _14282_/X VGND VGND VPWR VPWR _20504_/B sky130_fd_sc_hd__o21a_4
X_21481_ _17720_/X VGND VGND VPWR VPWR _21481_/X sky130_fd_sc_hd__buf_2
XFILLER_119_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14426__A _14408_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20432_ _20447_/A _20431_/Y VGND VGND VPWR VPWR _20451_/A sky130_fd_sc_hd__and2_4
X_23220_ _22545_/X _23219_/X _23044_/X _11753_/A _23111_/X VGND VGND VPWR VPWR _23220_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16307__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21300__B1 _24704_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22643__A _22611_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20363_ _23394_/Q VGND VGND VPWR VPWR _22234_/B sky130_fd_sc_hd__inv_2
X_23151_ _22654_/A VGND VGND VPWR VPWR _23310_/B sky130_fd_sc_hd__buf_2
Xclkbuf_5_0_0_HCLK clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_106_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22102_ _20699_/Y _21105_/A VGND VGND VPWR VPWR _22102_/X sky130_fd_sc_hd__or2_4
X_23082_ _24591_/Q _23082_/B VGND VGND VPWR VPWR _23082_/X sky130_fd_sc_hd__or2_4
X_20294_ _23420_/Q VGND VGND VPWR VPWR _20294_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22033_ _21681_/A _22012_/Y _22019_/Y _22026_/Y _22032_/Y VGND VGND VPWR VPWR _22033_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__11785__A _11777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22800__B1 _22797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22159__A2 _21352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23984_ _24322_/CLK _23983_/Q HRESETn VGND VGND VPWR VPWR _23984_/Q sky130_fd_sc_hd__dfrtp_4
X_22935_ _24654_/Q _22722_/B VGND VGND VPWR VPWR _22935_/X sky130_fd_sc_hd__or2_4
XFILLER_44_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15046__B1 _25022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_HCLK_A clkbuf_3_6_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22866_ _15791_/A _22865_/X _22485_/X _25525_/Q _22775_/X VGND VGND VPWR VPWR _22866_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22818__A _22270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24605_ _24600_/CLK _24605_/D HRESETn VGND VGND VPWR VPWR _22273_/A sky130_fd_sc_hd__dfrtp_4
X_21817_ _20329_/A _20318_/X _23383_/Q _21995_/A VGND VGND VPWR VPWR _21817_/X sky130_fd_sc_hd__o22a_4
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24103__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22797_ _22923_/A VGND VGND VPWR VPWR _22797_/X sky130_fd_sc_hd__buf_2
XFILLER_52_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16816__A _16807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12550_ _25397_/Q _24851_/Q _12708_/A _12549_/Y VGND VGND VPWR VPWR _12557_/B sky130_fd_sc_hd__o22a_4
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24536_ _24541_/CLK _24536_/D HRESETn VGND VGND VPWR VPWR _16535_/A sky130_fd_sc_hd__dfrtp_4
X_21748_ _21629_/A _21748_/B VGND VGND VPWR VPWR _21750_/B sky130_fd_sc_hd__or2_4
XANTENNA__16546__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16929__A2_N _16927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _12481_/A VGND VGND VPWR VPWR _12481_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24467_ _24033_/CLK _24467_/D HRESETn VGND VGND VPWR VPWR _16716_/A sky130_fd_sc_hd__dfrtp_4
X_21679_ _18291_/X VGND VGND VPWR VPWR _21679_/X sky130_fd_sc_hd__buf_2
XFILLER_138_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ _14220_/A VGND VGND VPWR VPWR _14221_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_16_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_16_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23418_ _23394_/CLK _23418_/D VGND VGND VPWR VPWR _23418_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_138_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25309__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24398_ _24398_/CLK _16869_/X HRESETn VGND VGND VPWR VPWR _20085_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_79_0_HCLK clkbuf_7_79_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_79_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14151_ _14129_/X _14150_/X _25125_/Q _14136_/X VGND VGND VPWR VPWR _14151_/Y sky130_fd_sc_hd__a22oi_4
X_23349_ VGND VGND VPWR VPWR _23349_/HI IRQ[15] sky130_fd_sc_hd__conb_1
XFILLER_137_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13102_ _13102_/A _13101_/Y VGND VGND VPWR VPWR _13103_/B sky130_fd_sc_hd__or2_4
XANTENNA__20748__A1_N _20743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14082_ _13977_/X _14081_/X _14078_/X _25221_/Q _14076_/X VGND VGND VPWR VPWR _14082_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12185__A1_N _12277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14324__A2 _23344_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22398__A2 _21095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13033_ _12299_/Y _13035_/B _13032_/Y VGND VGND VPWR VPWR _13033_/X sky130_fd_sc_hd__o21a_4
X_17910_ _17909_/Y _17905_/Y _17909_/A _17905_/A VGND VGND VPWR VPWR _17910_/X sky130_fd_sc_hd__o22a_4
X_25019_ _25020_/CLK _15201_/Y HRESETn VGND VGND VPWR VPWR _25019_/Q sky130_fd_sc_hd__dfrtp_4
X_18890_ _18869_/X _18883_/X _24107_/Q _24108_/Q _18886_/X VGND VGND VPWR VPWR _18890_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_3_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17841_ _17759_/A _17841_/B VGND VGND VPWR VPWR _17842_/C sky130_fd_sc_hd__or2_4
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14984_ _14951_/X _14984_/B _14984_/C _14983_/X VGND VGND VPWR VPWR _14984_/X sky130_fd_sc_hd__or4_4
X_17772_ _16916_/Y _16948_/X _17771_/X VGND VGND VPWR VPWR _17772_/X sky130_fd_sc_hd__or3_4
XFILLER_43_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19511_ _19511_/A VGND VGND VPWR VPWR _21181_/B sky130_fd_sc_hd__inv_2
XFILLER_75_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13935_ _13953_/A _13932_/Y _13924_/X _13935_/D VGND VGND VPWR VPWR _13936_/A sky130_fd_sc_hd__or4_4
X_16723_ _16723_/A VGND VGND VPWR VPWR _23021_/A sky130_fd_sc_hd__buf_2
XFILLER_78_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16654_ _16653_/Y _16651_/X _16386_/X _16651_/X VGND VGND VPWR VPWR _24493_/D sky130_fd_sc_hd__a2bb2o_4
X_19442_ _18204_/B VGND VGND VPWR VPWR _19442_/Y sky130_fd_sc_hd__inv_2
X_13866_ _20663_/A _13861_/X _22172_/A _13863_/X VGND VGND VPWR VPWR _13866_/X sky130_fd_sc_hd__o22a_4
X_15605_ _15588_/A VGND VGND VPWR VPWR _15605_/X sky130_fd_sc_hd__buf_2
X_12817_ _12886_/A _24794_/Q _12843_/A _12755_/Y VGND VGND VPWR VPWR _12817_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16585_ _16585_/A VGND VGND VPWR VPWR _16585_/Y sky130_fd_sc_hd__inv_2
X_19373_ _19372_/Y _19369_/X _19349_/X _19369_/X VGND VGND VPWR VPWR _19373_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22858__B1 _12555_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13797_ _16355_/A VGND VGND VPWR VPWR _13797_/X sky130_fd_sc_hd__buf_2
X_15536_ _12059_/X _15535_/X HADDR[4] _15535_/X VGND VGND VPWR VPWR _15536_/X sky130_fd_sc_hd__a2bb2o_4
X_18324_ _17465_/X _17451_/Y _17459_/X _19683_/B VGND VGND VPWR VPWR _18325_/A sky130_fd_sc_hd__and4_4
X_12748_ _25361_/Q _12746_/Y _12880_/A _23181_/A VGND VGND VPWR VPWR _12751_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18255_ _18235_/A _18253_/X _18254_/X _24216_/Q _18231_/A VGND VGND VPWR VPWR _18255_/X
+ sky130_fd_sc_hd__a32o_4
X_15467_ _15467_/A VGND VGND VPWR VPWR _15467_/Y sky130_fd_sc_hd__inv_2
X_12679_ _12679_/A _12689_/B VGND VGND VPWR VPWR _12686_/B sky130_fd_sc_hd__or2_4
XFILLER_129_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17206_ _17245_/C VGND VGND VPWR VPWR _17206_/X sky130_fd_sc_hd__buf_2
XFILLER_15_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14418_ _16528_/A VGND VGND VPWR VPWR _14418_/X sky130_fd_sc_hd__buf_2
X_18186_ _18186_/A _23830_/Q VGND VGND VPWR VPWR _18188_/B sky130_fd_sc_hd__or2_4
XANTENNA__23283__B1 _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15398_ _15301_/D _15398_/B VGND VGND VPWR VPWR _15398_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__20097__B1 _20096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17137_ _17041_/C _17135_/X _17136_/Y VGND VGND VPWR VPWR _17137_/X sky130_fd_sc_hd__o21a_4
X_14349_ _14338_/A _14348_/Y VGND VGND VPWR VPWR _14349_/X sky130_fd_sc_hd__or2_4
XANTENNA__17557__A _24701_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16461__A _16461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17068_ _17005_/Y _17066_/X _17067_/X _17061_/Y VGND VGND VPWR VPWR _17068_/X sky130_fd_sc_hd__a211o_4
X_16019_ _24725_/Q VGND VGND VPWR VPWR _16019_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15077__A _15077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24685__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17292__A _17257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21526__B _22879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24614__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19709_ _13247_/B VGND VGND VPWR VPWR _19709_/Y sky130_fd_sc_hd__inv_2
X_20981_ _22161_/A _23925_/Q _20982_/B VGND VGND VPWR VPWR _23924_/D sky130_fd_sc_hd__o21a_4
XFILLER_81_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0_0_HCLK_A clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22720_ _22520_/A VGND VGND VPWR VPWR _22796_/B sky130_fd_sc_hd__buf_2
XFILLER_80_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22651_ _22651_/A _23269_/B VGND VGND VPWR VPWR _22651_/X sky130_fd_sc_hd__or2_4
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21602_ _21595_/A VGND VGND VPWR VPWR _21629_/A sky130_fd_sc_hd__buf_2
X_25370_ _25368_/CLK _25370_/D HRESETn VGND VGND VPWR VPWR _12926_/A sky130_fd_sc_hd__dfrtp_4
X_22582_ _22581_/X VGND VGND VPWR VPWR _22582_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21521__B1 _12552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24321_ _24955_/CLK _17411_/X HRESETn VGND VGND VPWR VPWR _21000_/A sky130_fd_sc_hd__dfrtp_4
X_21533_ _21418_/X VGND VGND VPWR VPWR _21533_/X sky130_fd_sc_hd__buf_2
XANTENNA__25473__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15200__B1 _15199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24252_ _24252_/CLK _24252_/D HRESETn VGND VGND VPWR VPWR _24252_/Q sky130_fd_sc_hd__dfrtp_4
X_21464_ _21460_/A _21462_/X _21464_/C VGND VGND VPWR VPWR _21464_/X sky130_fd_sc_hd__and3_4
XANTENNA__15751__A1 _15749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25402__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23203_ _23133_/A _23203_/B _23203_/C VGND VGND VPWR VPWR _23203_/X sky130_fd_sc_hd__and3_4
X_20415_ _20414_/Y _20412_/X _18267_/X _20412_/X VGND VGND VPWR VPWR _23372_/D sky130_fd_sc_hd__a2bb2o_4
X_21395_ _21391_/X _21394_/X _21233_/X VGND VGND VPWR VPWR _21395_/X sky130_fd_sc_hd__o21a_4
X_24183_ _24373_/CLK _18378_/X HRESETn VGND VGND VPWR VPWR _24183_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16371__A _16371_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23134_ _24592_/Q _23171_/B VGND VGND VPWR VPWR _23137_/B sky130_fd_sc_hd__or2_4
X_20346_ _22013_/B _20340_/X _19618_/A _20345_/X VGND VGND VPWR VPWR _20346_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20277_ _20276_/X VGND VGND VPWR VPWR _20290_/A sky130_fd_sc_hd__inv_2
X_23065_ _23065_/A _23065_/B _23064_/X VGND VGND VPWR VPWR _23066_/D sky130_fd_sc_hd__and3_4
XFILLER_89_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22016_ _22016_/A _22016_/B VGND VGND VPWR VPWR _22016_/X sky130_fd_sc_hd__or2_4
XFILLER_103_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24355__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11981_ _11654_/A _11654_/B _11976_/X VGND VGND VPWR VPWR _11981_/X sky130_fd_sc_hd__and3_4
XFILLER_112_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21155__C _21314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23967_ _23967_/CLK _20995_/B HRESETn VGND VGND VPWR VPWR _14796_/C sky130_fd_sc_hd__dfstp_4
XFILLER_57_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13720_ _11663_/Y _13685_/X VGND VGND VPWR VPWR _13720_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__14227__A1_N _14226_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22918_ _23054_/A _22918_/B VGND VGND VPWR VPWR _22918_/Y sky130_fd_sc_hd__nor2_4
X_23898_ _23905_/CLK _18953_/X VGND VGND VPWR VPWR _18951_/A sky130_fd_sc_hd__dfxtp_4
X_13651_ _13651_/A VGND VGND VPWR VPWR _13653_/A sky130_fd_sc_hd__inv_2
XFILLER_71_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22849_ _22849_/A VGND VGND VPWR VPWR _22849_/Y sky130_fd_sc_hd__inv_2
X_12602_ _12602_/A VGND VGND VPWR VPWR _12664_/A sky130_fd_sc_hd__buf_2
XFILLER_13_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22267__B _22266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16370_ _16722_/A VGND VGND VPWR VPWR _22441_/A sky130_fd_sc_hd__buf_2
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A VGND VGND VPWR VPWR _13582_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16519__B1 _16147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15321_ _15320_/X VGND VGND VPWR VPWR _15322_/B sky130_fd_sc_hd__inv_2
XANTENNA__23990__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12533_ _12533_/A VGND VGND VPWR VPWR _12533_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24519_ _24553_/CLK _16580_/X HRESETn VGND VGND VPWR VPWR _24519_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25499_ _25497_/CLK _11918_/X HRESETn VGND VGND VPWR VPWR _25499_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18040_ _17928_/X _18040_/B _18040_/C VGND VGND VPWR VPWR _18040_/X sky130_fd_sc_hd__and3_4
X_15252_ _15252_/A VGND VGND VPWR VPWR _15253_/B sky130_fd_sc_hd__inv_2
XFILLER_9_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12464_ _12429_/X _12464_/B _12464_/C VGND VGND VPWR VPWR _25433_/D sky130_fd_sc_hd__and3_4
XANTENNA__25143__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22283__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14203_ _20506_/A VGND VGND VPWR VPWR _20500_/A sky130_fd_sc_hd__inv_2
XFILLER_138_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17377__A _17199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15183_ _15183_/A VGND VGND VPWR VPWR _25023_/D sky130_fd_sc_hd__inv_2
X_12395_ _12266_/Y _12392_/X _12387_/B _12394_/X VGND VGND VPWR VPWR _12396_/A sky130_fd_sc_hd__a211o_4
XANTENNA__17808__C _17792_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14134_ _23949_/D _14133_/X _14416_/A _23949_/D VGND VGND VPWR VPWR _25210_/D sky130_fd_sc_hd__a2bb2o_4
X_19991_ _19991_/A VGND VGND VPWR VPWR _19991_/X sky130_fd_sc_hd__buf_2
XFILLER_10_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_103_0_HCLK clkbuf_7_51_0_HCLK/X VGND VGND VPWR VPWR _24643_/CLK sky130_fd_sc_hd__clkbuf_1
X_14065_ _14081_/A VGND VGND VPWR VPWR _14065_/X sky130_fd_sc_hd__buf_2
X_18942_ _23901_/Q VGND VGND VPWR VPWR _18942_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_166_0_HCLK clkbuf_7_83_0_HCLK/X VGND VGND VPWR VPWR _23623_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_9_0_HCLK clkbuf_7_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13016_ _13038_/A _13014_/X _13015_/X VGND VGND VPWR VPWR _25351_/D sky130_fd_sc_hd__and3_4
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18873_ _18873_/A _18873_/B VGND VGND VPWR VPWR _18874_/B sky130_fd_sc_hd__or2_4
XFILLER_94_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22791__A2 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17824_ _17834_/A _17824_/B _17823_/Y VGND VGND VPWR VPWR _17824_/X sky130_fd_sc_hd__and3_4
XANTENNA__15625__A _15625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24096__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11819__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14967_ _24429_/Q VGND VGND VPWR VPWR _14967_/Y sky130_fd_sc_hd__inv_2
X_17755_ _24259_/Q VGND VGND VPWR VPWR _17755_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24025__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13145__A _13233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16706_ _24471_/Q VGND VGND VPWR VPWR _16706_/Y sky130_fd_sc_hd__inv_2
X_13918_ _13918_/A _13897_/X _13918_/C _13918_/D VGND VGND VPWR VPWR _13965_/B sky130_fd_sc_hd__and4_4
X_14898_ _15067_/D VGND VGND VPWR VPWR _15219_/C sky130_fd_sc_hd__buf_2
X_17686_ _17576_/Y _17662_/X _17683_/Y _17601_/X VGND VGND VPWR VPWR _17686_/X sky130_fd_sc_hd__a211o_4
XFILLER_90_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21751__B1 _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22458__A _22783_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19425_ _19431_/A VGND VGND VPWR VPWR _19425_/X sky130_fd_sc_hd__buf_2
X_13849_ _13848_/Y _13822_/A _13810_/X _13822_/A VGND VGND VPWR VPWR _25242_/D sky130_fd_sc_hd__a2bb2o_4
X_16637_ _16637_/A VGND VGND VPWR VPWR _24499_/D sky130_fd_sc_hd__inv_2
XFILLER_35_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19356_ _19355_/Y VGND VGND VPWR VPWR _19356_/X sky130_fd_sc_hd__buf_2
XFILLER_50_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16568_ _16567_/Y _16563_/X _16398_/X _16563_/X VGND VGND VPWR VPWR _16568_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14784__A2 _16880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18307_ _21173_/A VGND VGND VPWR VPWR _18307_/X sky130_fd_sc_hd__buf_2
X_15519_ _11730_/A VGND VGND VPWR VPWR _15519_/Y sky130_fd_sc_hd__inv_2
X_16499_ _16504_/A VGND VGND VPWR VPWR _16499_/X sky130_fd_sc_hd__buf_2
X_19287_ _19287_/A VGND VGND VPWR VPWR _19287_/Y sky130_fd_sc_hd__inv_2
X_18238_ _18231_/A VGND VGND VPWR VPWR _18238_/X sky130_fd_sc_hd__buf_2
XFILLER_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20706__A _20678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12547__B2 _12546_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18169_ _18201_/A _18169_/B _18169_/C VGND VGND VPWR VPWR _18170_/C sky130_fd_sc_hd__and3_4
XFILLER_11_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16191__A _23242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14704__A _14675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16931__A1_N _16130_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_62_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20200_ _20200_/A VGND VGND VPWR VPWR _21749_/B sky130_fd_sc_hd__inv_2
X_21180_ _24202_/Q _21171_/X _21180_/C VGND VGND VPWR VPWR _21180_/X sky130_fd_sc_hd__or3_4
XANTENNA__24866__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15497__B1 HADDR[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20131_ _22192_/B _20128_/X _20082_/X _20128_/X VGND VGND VPWR VPWR _23483_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12224__A _21526_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20062_ _20061_/Y _20057_/X _19841_/X _20057_/A VGND VGND VPWR VPWR _20062_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15535__A _15535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24870_ _24852_/CLK _24870_/D HRESETn VGND VGND VPWR VPWR _24870_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16997__B1 _16039_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22519__C1 _22518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23821_ _25044_/CLK _19172_/X VGND VGND VPWR VPWR _18219_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_22_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23752_ _23772_/CLK _23752_/D VGND VGND VPWR VPWR _23752_/Q sky130_fd_sc_hd__dfxtp_4
X_20964_ _12130_/X _20965_/B VGND VGND VPWR VPWR _20964_/X sky130_fd_sc_hd__and2_4
XANTENNA__22368__A _21618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17410__A1 _17387_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22703_ _22703_/A _21511_/X _21859_/C VGND VGND VPWR VPWR _22703_/X sky130_fd_sc_hd__and3_4
XFILLER_53_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17410__B2 _17404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23683_ _23683_/CLK _19565_/X VGND VGND VPWR VPWR _23683_/Q sky130_fd_sc_hd__dfxtp_4
X_20895_ _20882_/X _20894_/Y _24483_/Q _20886_/X VGND VGND VPWR VPWR _20895_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25422_ _25368_/CLK _25422_/D HRESETn VGND VGND VPWR VPWR _25422_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22634_ _22634_/A _22598_/B VGND VGND VPWR VPWR _22634_/X sky130_fd_sc_hd__and2_4
XANTENNA__16085__B _22493_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12786__A1 _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25353_ _23370_/CLK _13006_/X HRESETn VGND VGND VPWR VPWR _25353_/Q sky130_fd_sc_hd__dfrtp_4
X_22565_ _21009_/X VGND VGND VPWR VPWR _22565_/X sky130_fd_sc_hd__buf_2
XANTENNA__22815__B _21048_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24304_ _25436_/CLK _17610_/Y HRESETn VGND VGND VPWR VPWR _24304_/Q sky130_fd_sc_hd__dfrtp_4
X_21516_ _23314_/B _21516_/B VGND VGND VPWR VPWR _21516_/X sky130_fd_sc_hd__and2_4
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15724__A1 _15548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25284_ _25284_/CLK _13675_/X HRESETn VGND VGND VPWR VPWR _23343_/B sky130_fd_sc_hd__dfrtp_4
X_22496_ _16599_/Y _22442_/X _21573_/X _22495_/X VGND VGND VPWR VPWR _22496_/X sky130_fd_sc_hd__o22a_4
X_24235_ _23828_/CLK _24235_/D HRESETn VGND VGND VPWR VPWR _24235_/Q sky130_fd_sc_hd__dfrtp_4
X_21447_ _21192_/A VGND VGND VPWR VPWR _21455_/A sky130_fd_sc_hd__buf_2
XANTENNA__18269__A3 _16270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25128__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12180_ _12179_/Y _24766_/Q _12179_/Y _24766_/Q VGND VGND VPWR VPWR _12186_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24166_ _24159_/CLK _24166_/D HRESETn VGND VGND VPWR VPWR _18400_/A sky130_fd_sc_hd__dfrtp_4
X_21378_ _21374_/X _21377_/X _21233_/X VGND VGND VPWR VPWR _21388_/B sky130_fd_sc_hd__o21a_4
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11854__A1_N _11850_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23117_ _23115_/X _23116_/X _23117_/C VGND VGND VPWR VPWR _23117_/X sky130_fd_sc_hd__or3_4
X_20329_ _20329_/A VGND VGND VPWR VPWR _21977_/B sky130_fd_sc_hd__buf_2
XFILLER_134_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24097_ _24097_/CLK _24097_/D HRESETn VGND VGND VPWR VPWR _24097_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17536__A2_N _17565_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24536__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22550__B _22590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_239_0_HCLK clkbuf_8_239_0_HCLK/A VGND VGND VPWR VPWR _25351_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_110_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21447__A _21192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23048_ _12244_/Y _22980_/X _24268_/Q _22906_/X VGND VGND VPWR VPWR _23048_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15870_ _12782_/Y _15869_/X _11749_/X _15869_/X VGND VGND VPWR VPWR _15870_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14821_ _25188_/Q _14810_/X _14811_/X _14820_/Y VGND VGND VPWR VPWR _14821_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24999_ _25002_/CLK _24999_/D HRESETn VGND VGND VPWR VPWR _14966_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_45_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19926__B1 _19797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14752_ _14752_/A _14744_/X VGND VGND VPWR VPWR _14752_/X sky130_fd_sc_hd__and2_4
X_17540_ _11844_/Y _17576_/A _11753_/A _17559_/A VGND VGND VPWR VPWR _17540_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ _11963_/X VGND VGND VPWR VPWR _11964_/X sky130_fd_sc_hd__buf_2
XANTENNA__22278__A _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13703_ _13713_/A VGND VGND VPWR VPWR _13703_/X sky130_fd_sc_hd__buf_2
X_17471_ _17489_/B VGND VGND VPWR VPWR _17471_/Y sky130_fd_sc_hd__inv_2
X_14683_ _14676_/X _14750_/A VGND VGND VPWR VPWR _14684_/A sky130_fd_sc_hd__and2_4
X_11895_ _25505_/Q _11893_/Y _11887_/X _11894_/X VGND VGND VPWR VPWR _25505_/D sky130_fd_sc_hd__o22a_4
XFILLER_72_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16276__A _22671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25395__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19210_ _19210_/A VGND VGND VPWR VPWR _19210_/Y sky130_fd_sc_hd__inv_2
X_13634_ _13634_/A VGND VGND VPWR VPWR _13635_/A sky130_fd_sc_hd__inv_2
X_16422_ _16421_/Y _16419_/X _16235_/X _16419_/X VGND VGND VPWR VPWR _16422_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25324__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16353_ _16352_/Y _16350_/X _16064_/X _16350_/X VGND VGND VPWR VPWR _16353_/X sky130_fd_sc_hd__a2bb2o_4
X_19141_ _18122_/B VGND VGND VPWR VPWR _19141_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13565_ _13565_/A VGND VGND VPWR VPWR _13565_/Y sky130_fd_sc_hd__inv_2
X_15304_ _15299_/X _15301_/X _15303_/X VGND VGND VPWR VPWR _15305_/C sky130_fd_sc_hd__or3_4
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12516_ _12595_/A _12514_/Y _12645_/A _12527_/A VGND VGND VPWR VPWR _12516_/X sky130_fd_sc_hd__a2bb2o_4
X_19072_ _19070_/Y _19068_/X _19071_/X _19068_/X VGND VGND VPWR VPWR _19072_/X sky130_fd_sc_hd__a2bb2o_4
X_16284_ _24629_/Q VGND VGND VPWR VPWR _16284_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15715__A1 _15548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23238__B1 _22797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13496_ _13533_/D _13496_/B _12066_/X _13495_/X VGND VGND VPWR VPWR _13497_/A sky130_fd_sc_hd__or4_4
XFILLER_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15235_ _15216_/A _15235_/B _15234_/X VGND VGND VPWR VPWR _25010_/D sky130_fd_sc_hd__and3_4
X_18023_ _14645_/A VGND VGND VPWR VPWR _18023_/X sky130_fd_sc_hd__buf_2
XFILLER_60_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12447_ _12447_/A VGND VGND VPWR VPWR _12448_/B sky130_fd_sc_hd__inv_2
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_49_0_HCLK clkbuf_6_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_99_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15166_ _15180_/A _15166_/B _15166_/C _15165_/X VGND VGND VPWR VPWR _15169_/B sky130_fd_sc_hd__or4_4
XANTENNA__18665__B1 _16616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20067__A3 _13835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12378_ _12378_/A VGND VGND VPWR VPWR _12993_/A sky130_fd_sc_hd__buf_2
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15479__B1 _14470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14117_ _14117_/A _14117_/B _14117_/C VGND VGND VPWR VPWR _14117_/X sky130_fd_sc_hd__or3_4
XFILLER_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15097_ _24982_/Q _15096_/A _15296_/A _15096_/Y VGND VGND VPWR VPWR _15097_/X sky130_fd_sc_hd__o22a_4
X_19974_ _19991_/A VGND VGND VPWR VPWR _19974_/X sky130_fd_sc_hd__buf_2
XFILLER_45_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24277__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14151__B1 _25125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14048_ _14009_/B VGND VGND VPWR VPWR _14049_/D sky130_fd_sc_hd__inv_2
X_18925_ _18937_/A VGND VGND VPWR VPWR _18925_/X sky130_fd_sc_hd__buf_2
XANTENNA__18417__B1 _16246_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21357__A _21139_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24206__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18856_ _24558_/Q _18675_/X _24558_/Q _18675_/X VGND VGND VPWR VPWR _18859_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20775__B2 _20774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17807_ _17737_/X VGND VGND VPWR VPWR _17834_/A sky130_fd_sc_hd__buf_2
Xclkbuf_4_4_0_HCLK clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18787_ _18792_/A _18792_/B _18608_/X _18792_/C VGND VGND VPWR VPWR _18788_/A sky130_fd_sc_hd__or4_4
XFILLER_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15999_ _24733_/Q VGND VGND VPWR VPWR _15999_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19917__B1 _19783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17738_ _17737_/X VGND VGND VPWR VPWR _17738_/X sky130_fd_sc_hd__buf_2
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23291__B _22832_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17669_ _17499_/Y _17672_/B VGND VGND VPWR VPWR _17673_/B sky130_fd_sc_hd__or2_4
X_19408_ _19401_/A VGND VGND VPWR VPWR _19408_/X sky130_fd_sc_hd__buf_2
XFILLER_126_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20680_ _20770_/A VGND VGND VPWR VPWR _20680_/X sky130_fd_sc_hd__buf_2
XFILLER_51_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25065__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21820__A _13784_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19339_ _19333_/Y VGND VGND VPWR VPWR _19339_/X sky130_fd_sc_hd__buf_2
XFILLER_108_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22350_ _17706_/A _22346_/X _22347_/X _22348_/X _22349_/X VGND VGND VPWR VPWR _22350_/X
+ sky130_fd_sc_hd__a32o_4
X_21301_ _22705_/A _21300_/X VGND VGND VPWR VPWR _21301_/X sky130_fd_sc_hd__and2_4
XFILLER_136_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13717__B1 _13714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22281_ _22281_/A _21858_/X VGND VGND VPWR VPWR _22281_/X sky130_fd_sc_hd__and2_4
XFILLER_129_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14434__A _21352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24020_ _24018_/CLK _20782_/Y HRESETn VGND VGND VPWR VPWR _20779_/A sky130_fd_sc_hd__dfrtp_4
X_21232_ _21250_/A _21229_/X _21231_/X VGND VGND VPWR VPWR _21232_/X sky130_fd_sc_hd__and3_4
XANTENNA__22452__A1 _12104_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13193__B2 _11970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21163_ _24199_/Q _21163_/B VGND VGND VPWR VPWR _21163_/X sky130_fd_sc_hd__or2_4
XFILLER_116_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20114_ _21892_/B _20111_/X _20089_/X _20111_/X VGND VGND VPWR VPWR _23489_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18408__B1 _16249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21267__A _13598_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21094_ _16075_/A _21049_/X _22962_/A _21093_/X VGND VGND VPWR VPWR _21094_/X sky130_fd_sc_hd__a211o_4
XFILLER_63_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20215__B1 _19755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15890__B1 _24787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20045_ _20057_/A VGND VGND VPWR VPWR _20045_/X sky130_fd_sc_hd__buf_2
X_24922_ _24923_/CLK _24922_/D HRESETn VGND VGND VPWR VPWR _11730_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_24_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_69_0_HCLK clkbuf_8_69_0_HCLK/A VGND VGND VPWR VPWR _24322_/CLK sky130_fd_sc_hd__clkbuf_1
X_24853_ _24018_/CLK _15753_/X HRESETn VGND VGND VPWR VPWR _24853_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17480__A _24310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23804_ _23660_/CLK _19223_/X VGND VGND VPWR VPWR _13182_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21714__B _21548_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24784_ _24800_/CLK _15893_/X HRESETn VGND VGND VPWR VPWR _22623_/A sky130_fd_sc_hd__dfrtp_4
X_21996_ _21996_/A _13817_/A VGND VGND VPWR VPWR _22384_/A sky130_fd_sc_hd__or2_4
XFILLER_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _23722_/CLK _19416_/X VGND VGND VPWR VPWR _18139_/B sky130_fd_sc_hd__dfxtp_4
X_20947_ _20943_/X VGND VGND VPWR VPWR _20947_/Y sky130_fd_sc_hd__inv_2
XPHY_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__B1 _12277_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _24223_/Q VGND VGND VPWR VPWR _22532_/A sky130_fd_sc_hd__inv_2
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23666_ _23545_/CLK _19620_/X VGND VGND VPWR VPWR _19617_/A sky130_fd_sc_hd__dfxtp_4
X_20878_ _20879_/B VGND VGND VPWR VPWR _20878_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22826__A _23069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25405_ _25400_/CLK _25405_/D HRESETn VGND VGND VPWR VPWR _25405_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21730__A _22923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22617_ _22511_/B _22614_/X _22413_/X _22616_/X VGND VGND VPWR VPWR _22617_/X sky130_fd_sc_hd__o22a_4
XFILLER_35_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22140__B1 _21024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23597_ _23598_/CLK _19820_/X VGND VGND VPWR VPWR _13459_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13350_ _13314_/A _13350_/B _13350_/C VGND VGND VPWR VPWR _13351_/C sky130_fd_sc_hd__or3_4
XFILLER_122_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25336_ _24852_/CLK _13069_/Y HRESETn VGND VGND VPWR VPWR _12349_/A sky130_fd_sc_hd__dfrtp_4
X_22548_ _22545_/X _22546_/X _22127_/C _24852_/Q _22547_/X VGND VGND VPWR VPWR _22549_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22691__B2 _22442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12301_ _12293_/X _12295_/X _12298_/X _12300_/X VGND VGND VPWR VPWR _12301_/X sky130_fd_sc_hd__or4_4
XANTENNA__24788__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13281_ _13156_/X VGND VGND VPWR VPWR _13421_/A sky130_fd_sc_hd__buf_2
X_25267_ _25055_/CLK _13756_/Y HRESETn VGND VGND VPWR VPWR _25267_/Q sky130_fd_sc_hd__dfrtp_4
X_22479_ _21295_/X VGND VGND VPWR VPWR _22479_/X sky130_fd_sc_hd__buf_2
X_15020_ _15241_/A _24446_/Q _15209_/A _15019_/Y VGND VGND VPWR VPWR _15021_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24717__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12232_ _22141_/A VGND VGND VPWR VPWR _12232_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24218_ _24214_/CLK _24218_/D HRESETn VGND VGND VPWR VPWR _11677_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_120_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22443__B2 _22442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25198_ _25098_/CLK _25198_/D HRESETn VGND VGND VPWR VPWR _14173_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_5_3_0_HCLK_A clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12163_ _12163_/A _12163_/B VGND VGND VPWR VPWR _12163_/X sky130_fd_sc_hd__and2_4
X_24149_ _24159_/CLK _18584_/Y HRESETn VGND VGND VPWR VPWR _24149_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24370__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12094_ _12093_/X VGND VGND VPWR VPWR _13533_/D sky130_fd_sc_hd__buf_2
X_16971_ _16964_/X _16966_/X _16971_/C _16971_/D VGND VGND VPWR VPWR _16971_/X sky130_fd_sc_hd__or4_4
XFILLER_111_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15479__A1_N _14876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12799__A _12799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18710_ _18705_/B _18697_/X VGND VGND VPWR VPWR _18711_/A sky130_fd_sc_hd__or2_4
XANTENNA__15881__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15922_ _15685_/X _15920_/Y _15677_/X _15920_/Y VGND VGND VPWR VPWR _15922_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19072__B1 _19071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19690_ _19697_/A VGND VGND VPWR VPWR _19690_/X sky130_fd_sc_hd__buf_2
X_18641_ _18680_/B VGND VGND VPWR VPWR _18786_/C sky130_fd_sc_hd__buf_2
X_15853_ _15852_/Y VGND VGND VPWR VPWR _22835_/A sky130_fd_sc_hd__buf_2
XFILLER_64_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15633__B1 _15474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15325__D _15316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14804_ _14804_/A VGND VGND VPWR VPWR _14806_/B sky130_fd_sc_hd__inv_2
X_18572_ _18555_/A _18572_/B _18571_/Y VGND VGND VPWR VPWR _24154_/D sky130_fd_sc_hd__and3_4
X_12996_ _12991_/X _12993_/X _12995_/X VGND VGND VPWR VPWR _13071_/B sky130_fd_sc_hd__or3_4
X_15784_ _15642_/A _15784_/B VGND VGND VPWR VPWR _15931_/A sky130_fd_sc_hd__or2_4
XANTENNA__25505__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17523_ _17516_/X _17518_/X _17520_/X _17522_/X VGND VGND VPWR VPWR _17523_/X sky130_fd_sc_hd__or4_4
X_11947_ _11947_/A VGND VGND VPWR VPWR _11947_/X sky130_fd_sc_hd__buf_2
X_14735_ _14734_/Y _14708_/X _25055_/Q _14707_/A VGND VGND VPWR VPWR _14736_/A sky130_fd_sc_hd__o22a_4
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14666_ _19038_/A _14659_/X _14665_/X VGND VGND VPWR VPWR _14666_/Y sky130_fd_sc_hd__a21oi_4
X_17454_ _24197_/Q VGND VGND VPWR VPWR _20231_/C sky130_fd_sc_hd__inv_2
X_11878_ _11878_/A _11878_/B VGND VGND VPWR VPWR _11879_/B sky130_fd_sc_hd__nand2_4
XFILLER_127_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13617_ _25059_/Q VGND VGND VPWR VPWR _13617_/Y sky130_fd_sc_hd__inv_2
X_16405_ HWDATA[19] VGND VGND VPWR VPWR _16405_/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_12_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_12_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_14597_ _14567_/B _14586_/X _14596_/Y _14590_/X _14559_/A VGND VGND VPWR VPWR _25077_/D
+ sky130_fd_sc_hd__a32o_4
X_17385_ _17344_/A _17347_/B _17384_/X VGND VGND VPWR VPWR _24328_/D sky130_fd_sc_hd__and3_4
X_19124_ _19124_/A VGND VGND VPWR VPWR _19124_/Y sky130_fd_sc_hd__inv_2
X_13548_ _25076_/Q VGND VGND VPWR VPWR _14598_/A sky130_fd_sc_hd__inv_2
X_16336_ _16336_/A VGND VGND VPWR VPWR _16336_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22682__B2 _22271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16453__B _16453_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16267_ _16265_/Y _16187_/A _16266_/X _16187_/A VGND VGND VPWR VPWR _24635_/D sky130_fd_sc_hd__a2bb2o_4
X_19055_ HWDATA[1] VGND VGND VPWR VPWR _19055_/X sky130_fd_sc_hd__buf_2
X_13479_ _25310_/Q VGND VGND VPWR VPWR _13479_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24458__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15218_ _15218_/A VGND VGND VPWR VPWR _25015_/D sky130_fd_sc_hd__inv_2
X_18006_ _18006_/A _18006_/B _18006_/C VGND VGND VPWR VPWR _18006_/X sky130_fd_sc_hd__or3_4
X_16198_ _16197_/Y _16193_/X _15944_/X _16193_/X VGND VGND VPWR VPWR _16198_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22471__A _23035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15149_ _24589_/Q VGND VGND VPWR VPWR _15149_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17565__A _17565_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19957_ _19964_/A VGND VGND VPWR VPWR _19957_/X sky130_fd_sc_hd__buf_2
XFILLER_87_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24040__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_222_0_HCLK clkbuf_8_223_0_HCLK/A VGND VGND VPWR VPWR _24462_/CLK sky130_fd_sc_hd__clkbuf_1
X_18908_ _22062_/B _18902_/X _16872_/X _18907_/X VGND VGND VPWR VPWR _23914_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19888_ _18275_/X _18278_/D _19888_/C VGND VGND VPWR VPWR _19889_/A sky130_fd_sc_hd__or3_4
XANTENNA__12502__A _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20748__B2 _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18839_ _24543_/Q _18630_/A _16515_/Y _18792_/A VGND VGND VPWR VPWR _18839_/X sky130_fd_sc_hd__o22a_4
XFILLER_3_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15624__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21850_ _24332_/Q _21220_/A VGND VGND VPWR VPWR _21854_/B sky130_fd_sc_hd__or2_4
XANTENNA__25246__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20801_ _20799_/A _13136_/X _20800_/X VGND VGND VPWR VPWR _20801_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_93_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21781_ _21781_/A _21504_/B VGND VGND VPWR VPWR _21781_/X sky130_fd_sc_hd__and2_4
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23520_ _24923_/CLK _20034_/X VGND VGND VPWR VPWR _20033_/A sky130_fd_sc_hd__dfxtp_4
X_20732_ _13132_/A _13132_/B _20731_/Y VGND VGND VPWR VPWR _20732_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23451_ _23798_/CLK _23451_/D VGND VGND VPWR VPWR _23451_/Q sky130_fd_sc_hd__dfxtp_4
X_20663_ _20663_/A _14282_/X VGND VGND VPWR VPWR _20665_/B sky130_fd_sc_hd__or2_4
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22122__B1 _24847_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22402_ _22402_/A _22266_/X VGND VGND VPWR VPWR _22402_/X sky130_fd_sc_hd__or2_4
XFILLER_136_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23382_ _24219_/CLK _23382_/D VGND VGND VPWR VPWR _23382_/Q sky130_fd_sc_hd__dfxtp_4
X_20594_ _20447_/A VGND VGND VPWR VPWR _20594_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24881__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20684__B1 _20680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25121_ _25113_/CLK _14445_/X HRESETn VGND VGND VPWR VPWR _25121_/Q sky130_fd_sc_hd__dfstp_4
X_22333_ _21942_/A _22333_/B VGND VGND VPWR VPWR _22333_/X sky130_fd_sc_hd__or2_4
XANTENNA__11788__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24199__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24810__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25052_ _25054_/CLK _14743_/X HRESETn VGND VGND VPWR VPWR _22038_/A sky130_fd_sc_hd__dfrtp_4
X_22264_ _21275_/X VGND VGND VPWR VPWR _22658_/A sky130_fd_sc_hd__buf_2
XFILLER_121_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24128__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24003_ _24035_/CLK _20705_/Y HRESETn VGND VGND VPWR VPWR _13128_/A sky130_fd_sc_hd__dfrtp_4
X_21215_ _21008_/B _15649_/A _15655_/A _20812_/A _15658_/A VGND VGND VPWR VPWR _21215_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_2_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22812__C _22812_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17475__A _17474_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_32_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_32_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22195_ _21238_/X _22192_/X _22194_/X VGND VGND VPWR VPWR _22195_/X sky130_fd_sc_hd__and3_4
XANTENNA__21709__B _22111_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21146_ _21139_/X _21141_/X _21144_/X _21145_/X VGND VGND VPWR VPWR _21146_/X sky130_fd_sc_hd__and4_4
X_21077_ _21030_/X _21076_/Y _24767_/Q _21030_/X VGND VGND VPWR VPWR _21077_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20028_ _20028_/A VGND VGND VPWR VPWR _22010_/B sky130_fd_sc_hd__inv_2
X_24905_ _24055_/CLK _15576_/X HRESETn VGND VGND VPWR VPWR _24905_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16819__A _16807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15615__B1 _11825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12850_ _12764_/Y _12850_/B _12850_/C _12753_/A VGND VGND VPWR VPWR _12851_/D sky130_fd_sc_hd__or4_4
XANTENNA__16132__A1_N _16130_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15723__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24836_ _24836_/CLK _15800_/X HRESETn VGND VGND VPWR VPWR _24836_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19517__A2_N _19516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11801_ _11798_/Y _11795_/X _11800_/X _11795_/X VGND VGND VPWR VPWR _25522_/D sky130_fd_sc_hd__a2bb2o_4
X_12781_ _12871_/A VGND VGND VPWR VPWR _12864_/A sky130_fd_sc_hd__inv_2
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24767_ _24806_/CLK _15929_/X HRESETn VGND VGND VPWR VPWR _24767_/Q sky130_fd_sc_hd__dfrtp_4
X_21979_ _21975_/Y _21976_/X _21977_/X _21978_/X VGND VGND VPWR VPWR _21979_/X sky130_fd_sc_hd__a211o_4
XFILLER_92_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14502_/X _14519_/X _25107_/Q _14517_/X VGND VGND VPWR VPWR _14520_/X sky130_fd_sc_hd__o22a_4
XPHY_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11732_ _11732_/A VGND VGND VPWR VPWR _21027_/A sky130_fd_sc_hd__buf_2
XPHY_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23718_ _23718_/CLK _19463_/X VGND VGND VPWR VPWR _19461_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__15918__A1 _13588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24698_ _24699_/CLK _16091_/X HRESETn VGND VGND VPWR VPWR _23278_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_42_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22556__A _22556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24969__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14451_ _14182_/Y _14448_/X _14400_/X _14436_/Y VGND VGND VPWR VPWR _14451_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11663_ _25274_/Q VGND VGND VPWR VPWR _11663_/Y sky130_fd_sc_hd__inv_2
XPHY_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23649_ _23649_/CLK _23649_/D VGND VGND VPWR VPWR _19671_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13402_/A _13402_/B VGND VGND VPWR VPWR _13403_/C sky130_fd_sc_hd__or2_4
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17170_ _22273_/A _17369_/A _16293_/Y _24355_/Q VGND VGND VPWR VPWR _17170_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14382_ _14394_/B _14380_/X _14383_/A VGND VGND VPWR VPWR _14382_/X sky130_fd_sc_hd__a21o_4
XFILLER_128_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16121_ _16120_/Y _16118_/X _15962_/X _16118_/X VGND VGND VPWR VPWR _16121_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_114_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_229_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13333_ _13366_/A _13333_/B _13332_/X VGND VGND VPWR VPWR _13333_/X sky130_fd_sc_hd__and3_4
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25319_ _25316_/CLK _25319_/D HRESETn VGND VGND VPWR VPWR _25319_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17540__B1 _11753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24551__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16052_ _16060_/A VGND VGND VPWR VPWR _16052_/X sky130_fd_sc_hd__buf_2
XANTENNA__22416__A1 _23281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13264_ _13260_/X _13261_/X _13263_/X VGND VGND VPWR VPWR _13264_/X sky130_fd_sc_hd__and3_4
X_15003_ _15003_/A VGND VGND VPWR VPWR _15003_/Y sky130_fd_sc_hd__inv_2
X_12215_ _12213_/A _22892_/A _12286_/C _12214_/Y VGND VGND VPWR VPWR _12215_/X sky130_fd_sc_hd__o22a_4
XFILLER_6_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13195_ _11984_/Y _13194_/Y _11976_/A VGND VGND VPWR VPWR _13195_/X sky130_fd_sc_hd__o21a_4
X_19811_ _19810_/Y _19808_/X _19715_/X _19808_/X VGND VGND VPWR VPWR _19811_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12146_ _12106_/Y _12130_/X _12131_/Y _12145_/X VGND VGND VPWR VPWR _12157_/A sky130_fd_sc_hd__a211o_4
XFILLER_116_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19742_ _13392_/B VGND VGND VPWR VPWR _19742_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13418__A _13450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12077_ _12076_/Y _12074_/X _11838_/X _12074_/X VGND VGND VPWR VPWR _25472_/D sky130_fd_sc_hd__a2bb2o_4
X_16954_ _16953_/X VGND VGND VPWR VPWR _17805_/A sky130_fd_sc_hd__inv_2
XFILLER_133_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15905_ _12796_/Y _15904_/X _15627_/X _15904_/X VGND VGND VPWR VPWR _24777_/D sky130_fd_sc_hd__a2bb2o_4
X_19673_ _19673_/A VGND VGND VPWR VPWR _19673_/Y sky130_fd_sc_hd__inv_2
X_16885_ _16879_/A VGND VGND VPWR VPWR _16885_/X sky130_fd_sc_hd__buf_2
XANTENNA__16729__A _16733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15606__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18624_ _24509_/Q _18623_/A _16606_/Y _18623_/Y VGND VGND VPWR VPWR _18624_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_8_52_0_HCLK clkbuf_8_53_0_HCLK/A VGND VGND VPWR VPWR _24383_/CLK sky130_fd_sc_hd__clkbuf_1
X_15836_ _15766_/A VGND VGND VPWR VPWR _15836_/X sky130_fd_sc_hd__buf_2
XFILLER_65_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18555_ _18555_/A _18553_/X _18554_/X VGND VGND VPWR VPWR _18555_/X sky130_fd_sc_hd__and3_4
X_12979_ _12979_/A _12979_/B _12978_/X VGND VGND VPWR VPWR _12979_/X sky130_fd_sc_hd__and3_4
X_15767_ _15749_/X _15765_/X _15766_/X _24846_/Q _15711_/A VGND VGND VPWR VPWR _24846_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_18_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18556__C1 _18487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18944__A _18944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17506_ _24297_/Q VGND VGND VPWR VPWR _17567_/A sky130_fd_sc_hd__inv_2
X_14718_ _21633_/A _14717_/X _21633_/A _14717_/X VGND VGND VPWR VPWR _14718_/X sky130_fd_sc_hd__a2bb2o_4
X_18486_ _18521_/A VGND VGND VPWR VPWR _18821_/B sky130_fd_sc_hd__inv_2
X_15698_ _14620_/B _15694_/X VGND VGND VPWR VPWR _15698_/X sky130_fd_sc_hd__and2_4
XANTENNA__22466__A _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17437_ _17436_/Y _17432_/X _16720_/X _17432_/A VGND VGND VPWR VPWR _24313_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14649_ _25062_/Q VGND VGND VPWR VPWR _17975_/A sky130_fd_sc_hd__inv_2
XANTENNA__22104__B1 _20837_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24639__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17368_ _17349_/A _17370_/B _17367_/Y VGND VGND VPWR VPWR _24335_/D sky130_fd_sc_hd__o21a_4
XFILLER_105_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16183__B _22444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19107_ _19106_/Y VGND VGND VPWR VPWR _19107_/X sky130_fd_sc_hd__buf_2
X_16319_ _16318_/Y _16316_/X _15962_/X _16316_/X VGND VGND VPWR VPWR _24617_/D sky130_fd_sc_hd__a2bb2o_4
X_17299_ _17298_/X VGND VGND VPWR VPWR _17299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17531__B1 _11802_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24292__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19038_ _19038_/A _19038_/B _19038_/C _19038_/D VGND VGND VPWR VPWR _19038_/X sky130_fd_sc_hd__and4_4
XFILLER_133_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23080__A1 _21409_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_19_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_19_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_21000_ _21000_/A _21000_/B VGND VGND VPWR VPWR _21000_/Y sky130_fd_sc_hd__nor2_4
XFILLER_114_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25498__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12232__A _22141_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25427__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22951_ _14969_/A _22833_/X _22090_/X _22950_/X VGND VGND VPWR VPWR _22952_/C sky130_fd_sc_hd__a211o_4
XANTENNA__22591__B1 _24818_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21902_ _21898_/X _21901_/X _14712_/A VGND VGND VPWR VPWR _21902_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25080__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22882_ _16452_/A _22882_/B _22882_/C VGND VGND VPWR VPWR _22889_/C sky130_fd_sc_hd__and3_4
XFILLER_23_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23135__A2 _22998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24621_ _24330_/CLK _16309_/X HRESETn VGND VGND VPWR VPWR _23009_/A sky130_fd_sc_hd__dfrtp_4
X_21833_ _21830_/X _21833_/B _21832_/X VGND VGND VPWR VPWR _21833_/X sky130_fd_sc_hd__and3_4
XFILLER_70_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17492__A1_N _11815_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24552_ _24553_/CLK _16494_/X HRESETn VGND VGND VPWR VPWR _24552_/Q sky130_fd_sc_hd__dfrtp_4
X_21764_ _21616_/A _21764_/B VGND VGND VPWR VPWR _21766_/B sky130_fd_sc_hd__or2_4
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21280__A _21280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23503_ _24208_/CLK _23503_/D VGND VGND VPWR VPWR _23503_/Q sky130_fd_sc_hd__dfxtp_4
X_20715_ _15616_/Y _20698_/X _20706_/X _20714_/Y VGND VGND VPWR VPWR _20715_/X sky130_fd_sc_hd__o22a_4
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24483_ _24413_/CLK _16679_/X HRESETn VGND VGND VPWR VPWR _24483_/Q sky130_fd_sc_hd__dfrtp_4
X_21695_ _21512_/X _21694_/X _21514_/X _24845_/Q _21520_/X VGND VGND VPWR VPWR _21696_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_106_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23434_ _23434_/CLK _23434_/D VGND VGND VPWR VPWR _23434_/Q sky130_fd_sc_hd__dfxtp_4
X_20646_ _17396_/A _17396_/B VGND VGND VPWR VPWR _20646_/Y sky130_fd_sc_hd__nand2_4
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24309__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23365_ _21008_/X VGND VGND VPWR VPWR IRQ[11] sky130_fd_sc_hd__buf_2
X_20577_ _20577_/A VGND VGND VPWR VPWR _23940_/D sky130_fd_sc_hd__inv_2
XANTENNA__12407__A _25447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25104_ _25113_/CLK _14486_/X HRESETn VGND VGND VPWR VPWR _25104_/Q sky130_fd_sc_hd__dfrtp_4
X_22316_ _15461_/Y _22316_/B VGND VGND VPWR VPWR _22316_/Y sky130_fd_sc_hd__nor2_4
XFILLER_30_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23296_ _24463_/Q _22654_/X _23172_/X VGND VGND VPWR VPWR _23296_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14887__B2 _24412_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25035_ _24171_/CLK _14854_/X HRESETn VGND VGND VPWR VPWR _25035_/Q sky130_fd_sc_hd__dfrtp_4
X_22247_ _22247_/A _22247_/B _22246_/X VGND VGND VPWR VPWR _22248_/C sky130_fd_sc_hd__and3_4
XFILLER_69_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12898__B1 _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12000_ _25298_/Q VGND VGND VPWR VPWR _12000_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16089__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21082__B1 _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22178_ _22172_/X _22174_/Y _22176_/Y _22177_/X _21547_/Y VGND VGND VPWR VPWR _22178_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21129_ _13536_/A _12093_/X _13465_/Y _12093_/X VGND VGND VPWR VPWR _21129_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23944__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21455__A _21455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13951_ _13951_/A VGND VGND VPWR VPWR _13952_/D sky130_fd_sc_hd__inv_2
XFILLER_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16549__A _24531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12902_ _22660_/A _12799_/X _12600_/X _12847_/X VGND VGND VPWR VPWR _12902_/X sky130_fd_sc_hd__or4_4
Xclkbuf_7_39_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_79_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13882_ _21142_/A _13860_/X _23428_/Q _13855_/X VGND VGND VPWR VPWR _13882_/X sky130_fd_sc_hd__o22a_4
X_16670_ _24486_/Q VGND VGND VPWR VPWR _16670_/Y sky130_fd_sc_hd__inv_2
X_12833_ _25361_/Q VGND VGND VPWR VPWR _12833_/Y sky130_fd_sc_hd__inv_2
X_15621_ _22407_/A _15617_/X _15620_/X _15617_/X VGND VGND VPWR VPWR _24887_/D sky130_fd_sc_hd__a2bb2o_4
X_24819_ _24821_/CLK _24819_/D HRESETn VGND VGND VPWR VPWR _24819_/Q sky130_fd_sc_hd__dfrtp_4
X_18340_ _17456_/Y _18340_/B VGND VGND VPWR VPWR _18340_/X sky130_fd_sc_hd__or2_4
X_12764_ _25373_/Q VGND VGND VPWR VPWR _12764_/Y sky130_fd_sc_hd__inv_2
X_15552_ _15777_/A VGND VGND VPWR VPWR _15552_/Y sky130_fd_sc_hd__inv_2
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16013__B1 _11764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _11714_/Y VGND VGND VPWR VPWR _11716_/A sky130_fd_sc_hd__buf_2
X_14503_ _20441_/C _14503_/B VGND VGND VPWR VPWR _14503_/Y sky130_fd_sc_hd__nor2_4
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _24062_/Q VGND VGND VPWR VPWR _15484_/B sky130_fd_sc_hd__inv_2
X_18271_ _18270_/X VGND VGND VPWR VPWR _18272_/A sky130_fd_sc_hd__buf_2
X_12695_ _12695_/A VGND VGND VPWR VPWR _12695_/Y sky130_fd_sc_hd__inv_2
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24732__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _23008_/A VGND VGND VPWR VPWR _17222_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14434_ _21352_/A VGND VGND VPWR VPWR _22316_/B sky130_fd_sc_hd__buf_2
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ _14355_/X _14364_/X _12081_/A _14360_/X VGND VGND VPWR VPWR _25145_/D sky130_fd_sc_hd__o22a_4
X_17153_ _17153_/A VGND VGND VPWR VPWR _24364_/D sky130_fd_sc_hd__inv_2
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13316_ _13316_/A _19671_/A VGND VGND VPWR VPWR _13318_/B sky130_fd_sc_hd__or2_4
X_16104_ _16103_/Y _16101_/X _11764_/X _16101_/X VGND VGND VPWR VPWR _16104_/X sky130_fd_sc_hd__a2bb2o_4
X_17084_ _17077_/X VGND VGND VPWR VPWR _17088_/B sky130_fd_sc_hd__inv_2
X_14296_ _14296_/A _14296_/B VGND VGND VPWR VPWR _14301_/B sky130_fd_sc_hd__or2_4
XANTENNA__21860__A2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14878__A1 _14876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13247_ _13246_/X _13247_/B VGND VGND VPWR VPWR _13250_/B sky130_fd_sc_hd__or2_4
X_16035_ _16060_/A VGND VGND VPWR VPWR _16035_/X sky130_fd_sc_hd__buf_2
XANTENNA__18004__A _18046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13178_ _13177_/Y VGND VGND VPWR VPWR _13366_/A sky130_fd_sc_hd__buf_2
XFILLER_123_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15827__B1 _11822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12129_ _12147_/B VGND VGND VPWR VPWR _12129_/Y sky130_fd_sc_hd__inv_2
X_17986_ _18201_/A _17983_/X _17986_/C VGND VGND VPWR VPWR _17993_/B sky130_fd_sc_hd__and3_4
XANTENNA__25520__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19725_ _19725_/A VGND VGND VPWR VPWR _19725_/Y sky130_fd_sc_hd__inv_2
X_16937_ _16933_/X _16937_/B _16937_/C _16936_/X VGND VGND VPWR VPWR _16952_/B sky130_fd_sc_hd__or4_4
XFILLER_38_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16459__A _16728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19656_ _19655_/Y _19653_/X _19462_/X _19653_/X VGND VGND VPWR VPWR _19656_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16868_ _16880_/A VGND VGND VPWR VPWR _16868_/X sky130_fd_sc_hd__buf_2
XANTENNA__16252__B1 _16057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18607_ _24123_/Q VGND VGND VPWR VPWR _18607_/Y sky130_fd_sc_hd__inv_2
X_15819_ _15819_/A VGND VGND VPWR VPWR _15819_/X sky130_fd_sc_hd__buf_2
XFILLER_93_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19587_ _19587_/A VGND VGND VPWR VPWR _19587_/X sky130_fd_sc_hd__buf_2
X_16799_ _16799_/A VGND VGND VPWR VPWR _16799_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18538_ _18420_/Y _18541_/B VGND VGND VPWR VPWR _18538_/Y sky130_fd_sc_hd__nand2_4
XFILLER_94_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22876__B2 _21211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16004__B1 _15940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18469_ _18416_/Y _18469_/B _18411_/Y _18393_/Y VGND VGND VPWR VPWR _18476_/A sky130_fd_sc_hd__or4_4
XANTENNA__24473__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20500_ _20500_/A _14281_/X VGND VGND VPWR VPWR _20500_/X sky130_fd_sc_hd__and2_4
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21480_ _21485_/A _21480_/B _21480_/C VGND VGND VPWR VPWR _21480_/X sky130_fd_sc_hd__and3_4
XANTENNA__24402__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20431_ _14496_/X VGND VGND VPWR VPWR _20431_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17504__B1 _11864_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21300__A1 _21280_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23150_ _22186_/A VGND VGND VPWR VPWR _23150_/X sky130_fd_sc_hd__buf_2
X_20362_ _22346_/B _20361_/X _19612_/A _20361_/X VGND VGND VPWR VPWR _23395_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22101_ _22101_/A _22101_/B _22101_/C _22101_/D VGND VGND VPWR VPWR _22101_/X sky130_fd_sc_hd__or4_4
XFILLER_134_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15538__A _15535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23081_ _23081_/A VGND VGND VPWR VPWR _23081_/Y sky130_fd_sc_hd__inv_2
X_20293_ _20292_/Y _20290_/X _19995_/X _20290_/X VGND VGND VPWR VPWR _23421_/D sky130_fd_sc_hd__a2bb2o_4
X_22032_ _21481_/X _22031_/X _17728_/A VGND VGND VPWR VPWR _22032_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_103_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15818__B1 _24823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25230__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25261__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21275__A _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23983_ _24322_/CLK scl_i_S5 HRESETn VGND VGND VPWR VPWR _23983_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23193__C _22132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21706__C _21048_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22934_ _22905_/X _22912_/X _22918_/Y _22933_/X VGND VGND VPWR VPWR HRDATA[19] sky130_fd_sc_hd__a211o_4
XANTENNA__17191__C _17187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16243__B1 _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22865_ _22865_/A _22864_/X VGND VGND VPWR VPWR _22865_/X sky130_fd_sc_hd__or2_4
XFILLER_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21816_ _24198_/Q _21816_/B VGND VGND VPWR VPWR _21816_/X sky130_fd_sc_hd__or2_4
X_24604_ _24600_/CLK _16353_/X HRESETn VGND VGND VPWR VPWR _16352_/A sky130_fd_sc_hd__dfrtp_4
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22796_ _24583_/Q _22796_/B VGND VGND VPWR VPWR _22801_/B sky130_fd_sc_hd__or2_4
XFILLER_71_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24535_ _24502_/CLK _24535_/D HRESETn VGND VGND VPWR VPWR _24535_/Q sky130_fd_sc_hd__dfrtp_4
X_21747_ _21631_/A _21747_/B _21746_/X VGND VGND VPWR VPWR _21747_/X sky130_fd_sc_hd__and3_4
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12480_ _12203_/X _12471_/X VGND VGND VPWR VPWR _12481_/A sky130_fd_sc_hd__or2_4
XFILLER_106_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24466_ _24496_/CLK _16721_/X HRESETn VGND VGND VPWR VPWR _16719_/A sky130_fd_sc_hd__dfrtp_4
X_21678_ _21452_/A _21676_/X _21678_/C VGND VGND VPWR VPWR _21678_/X sky130_fd_sc_hd__and3_4
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22834__A _22923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24143__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23417_ _23714_/CLK _23417_/D VGND VGND VPWR VPWR _20303_/A sky130_fd_sc_hd__dfxtp_4
X_20629_ _20629_/A _20625_/A VGND VGND VPWR VPWR _20630_/B sky130_fd_sc_hd__nand2_4
XANTENNA__22095__A2 _21352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17928__A _17928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23292__A1 _24564_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24397_ _24396_/CLK _16873_/X HRESETn VGND VGND VPWR VPWR _20089_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_20_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22553__B _22592_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14150_ _25205_/Q _14101_/B _25205_/Q _14101_/B VGND VGND VPWR VPWR _14150_/X sky130_fd_sc_hd__a2bb2o_4
X_23348_ VGND VGND VPWR VPWR _23348_/HI IRQ[14] sky130_fd_sc_hd__conb_1
XFILLER_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13101_ _13081_/X VGND VGND VPWR VPWR _13101_/Y sky130_fd_sc_hd__inv_2
X_14081_ _14081_/A VGND VGND VPWR VPWR _14081_/X sky130_fd_sc_hd__buf_2
XANTENNA__19380__A2_N _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23279_ _22545_/X _23278_/X _22127_/C _25537_/Q _23111_/X VGND VGND VPWR VPWR _23279_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25349__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13032_ _12299_/Y _13035_/B _13031_/X VGND VGND VPWR VPWR _13032_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_65_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12335__A2 _24809_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25018_ _25020_/CLK _15204_/X HRESETn VGND VGND VPWR VPWR _25018_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17840_ _17752_/A _17840_/B VGND VGND VPWR VPWR _17840_/X sky130_fd_sc_hd__or2_4
XANTENNA__19581__C _13777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16482__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17771_ _17771_/A _17771_/B VGND VGND VPWR VPWR _17771_/X sky130_fd_sc_hd__or2_4
XFILLER_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14983_ _14976_/X _14978_/X _14979_/X _14982_/X VGND VGND VPWR VPWR _14983_/X sky130_fd_sc_hd__or4_4
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16279__A _22493_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21358__B2 _21548_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19510_ _19509_/Y _19507_/X _11955_/X _19507_/X VGND VGND VPWR VPWR _19510_/X sky130_fd_sc_hd__a2bb2o_4
X_16722_ _16722_/A VGND VGND VPWR VPWR _16723_/A sky130_fd_sc_hd__inv_2
X_13934_ _13957_/B _13956_/A _13889_/X _13930_/D VGND VGND VPWR VPWR _13935_/D sky130_fd_sc_hd__or4_4
XANTENNA__15037__B2 _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24984__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19441_ _19440_/Y _19438_/X _19349_/X _19438_/X VGND VGND VPWR VPWR _23726_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21913__A _17717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16653_ _16653_/A VGND VGND VPWR VPWR _16653_/Y sky130_fd_sc_hd__inv_2
X_13865_ _13852_/X _13864_/X VGND VGND VPWR VPWR _13865_/X sky130_fd_sc_hd__or2_4
XANTENNA__18494__A _18481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24913__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15604_ _15604_/A VGND VGND VPWR VPWR _15604_/Y sky130_fd_sc_hd__inv_2
X_12816_ _25377_/Q VGND VGND VPWR VPWR _12886_/A sky130_fd_sc_hd__inv_2
X_19372_ _18164_/B VGND VGND VPWR VPWR _19372_/Y sky130_fd_sc_hd__inv_2
X_16584_ _16581_/Y _16583_/X _16325_/X _16583_/X VGND VGND VPWR VPWR _16584_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13134__C _20761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13796_ _13795_/X VGND VGND VPWR VPWR _13796_/X sky130_fd_sc_hd__buf_2
XFILLER_50_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_126_0_HCLK clkbuf_7_63_0_HCLK/X VGND VGND VPWR VPWR _24572_/CLK sky130_fd_sc_hd__clkbuf_1
X_18323_ _24196_/Q VGND VGND VPWR VPWR _19683_/B sky130_fd_sc_hd__buf_2
X_15535_ _15535_/A VGND VGND VPWR VPWR _15535_/X sky130_fd_sc_hd__buf_2
X_12747_ _12747_/A VGND VGND VPWR VPWR _12880_/A sky130_fd_sc_hd__inv_2
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_189_0_HCLK clkbuf_7_94_0_HCLK/X VGND VGND VPWR VPWR _25425_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18254_ _18254_/A VGND VGND VPWR VPWR _18254_/X sky130_fd_sc_hd__buf_2
X_12678_ _12609_/A _12682_/B _12677_/Y VGND VGND VPWR VPWR _25407_/D sky130_fd_sc_hd__o21a_4
X_15466_ _15465_/Y _15463_/X _14414_/X _15463_/X VGND VGND VPWR VPWR _24944_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17205_ _24329_/Q VGND VGND VPWR VPWR _17245_/C sky130_fd_sc_hd__inv_2
XFILLER_54_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14417_ HWDATA[5] VGND VGND VPWR VPWR _16528_/A sky130_fd_sc_hd__buf_2
X_18185_ _18185_/A _18185_/B _18184_/X VGND VGND VPWR VPWR _18185_/X sky130_fd_sc_hd__or3_4
XANTENNA__22086__A2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15397_ _15073_/Y _15399_/B _15396_/Y VGND VGND VPWR VPWR _15397_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12047__A _16371_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17136_ _17041_/C _17135_/X _17056_/X VGND VGND VPWR VPWR _17136_/Y sky130_fd_sc_hd__a21oi_4
X_14348_ _14348_/A VGND VGND VPWR VPWR _14348_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11782__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16593__A1_N _16592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14279_ _14279_/A VGND VGND VPWR VPWR _15449_/A sky130_fd_sc_hd__buf_2
X_17067_ _17384_/B VGND VGND VPWR VPWR _17067_/X sky130_fd_sc_hd__buf_2
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16018_ _16017_/Y _16015_/X _11771_/X _16015_/X VGND VGND VPWR VPWR _16018_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25019__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21095__A _21306_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17969_ _18204_/A _17969_/B VGND VGND VPWR VPWR _17969_/X sky130_fd_sc_hd__or2_4
X_19708_ _19704_/Y _19707_/X _19664_/X _19707_/X VGND VGND VPWR VPWR _23636_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19411__B1 _19364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20980_ _23926_/Q VGND VGND VPWR VPWR _20982_/B sky130_fd_sc_hd__inv_2
XFILLER_66_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19639_ _19638_/Y VGND VGND VPWR VPWR _19639_/X sky130_fd_sc_hd__buf_2
XANTENNA__21823__A _21707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_22_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24654__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_85_0_HCLK clkbuf_7_85_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_85_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22650_ _22464_/A VGND VGND VPWR VPWR _23269_/B sky130_fd_sc_hd__buf_2
XANTENNA__21542__B _22111_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21601_ _21601_/A VGND VGND VPWR VPWR _21609_/A sky130_fd_sc_hd__buf_2
XFILLER_0_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22581_ _22511_/B _22578_/X _22413_/X _22580_/X VGND VGND VPWR VPWR _22581_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12245__A1_N _12244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21521__A1 _21512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21521__B2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16546__A1_N _16541_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24320_ _25192_/CLK _17419_/X HRESETn VGND VGND VPWR VPWR _20657_/A sky130_fd_sc_hd__dfrtp_4
X_21532_ _21295_/X VGND VGND VPWR VPWR _21532_/X sky130_fd_sc_hd__buf_2
XFILLER_138_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22654__A _22654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24251_ _24673_/CLK _24251_/D HRESETn VGND VGND VPWR VPWR _22181_/A sky130_fd_sc_hd__dfrtp_4
X_21463_ _21658_/A _20016_/Y VGND VGND VPWR VPWR _21464_/C sky130_fd_sc_hd__or2_4
XANTENNA__15751__A2 _15742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23202_ _24529_/Q _22467_/X _22834_/X _23201_/X VGND VGND VPWR VPWR _23203_/C sky130_fd_sc_hd__a211o_4
X_20414_ _23372_/Q VGND VGND VPWR VPWR _20414_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24182_ _24373_/CLK _18380_/X HRESETn VGND VGND VPWR VPWR _24182_/Q sky130_fd_sc_hd__dfrtp_4
X_21394_ _21398_/A _21392_/X _21394_/C VGND VGND VPWR VPWR _21394_/X sky130_fd_sc_hd__and3_4
XFILLER_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11796__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23133_ _23133_/A _23129_/X _23133_/C VGND VGND VPWR VPWR _23133_/X sky130_fd_sc_hd__and3_4
X_20345_ _20339_/Y VGND VGND VPWR VPWR _20345_/X sky130_fd_sc_hd__buf_2
XANTENNA__25442__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23064_ _24424_/Q _22929_/X _22997_/X _23063_/X VGND VGND VPWR VPWR _23064_/X sky130_fd_sc_hd__a211o_4
X_20276_ _20338_/A _19971_/X _20276_/C VGND VGND VPWR VPWR _20276_/X sky130_fd_sc_hd__or3_4
XFILLER_89_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22015_ _21671_/A _22015_/B _22014_/X VGND VGND VPWR VPWR _22015_/X sky130_fd_sc_hd__and3_4
XFILLER_130_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16464__B1 _16285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23329__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11980_ _11701_/A _11655_/A _11977_/X _11653_/A _11979_/X VGND VGND VPWR VPWR _11980_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19402__B1 _19313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23966_ _23964_/CLK _23966_/D HRESETn VGND VGND VPWR VPWR _23968_/D sky130_fd_sc_hd__dfstp_4
XFILLER_90_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22917_ _22783_/X _22914_/X _22786_/X _22916_/X VGND VGND VPWR VPWR _22918_/B sky130_fd_sc_hd__o22a_4
X_23897_ _23905_/CLK _18956_/X VGND VGND VPWR VPWR _13308_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16827__A _24416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24395__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13650_ _24050_/Q _24049_/Q _24051_/Q _20900_/B VGND VGND VPWR VPWR _13650_/X sky130_fd_sc_hd__or4_4
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22848_ _22753_/X _22845_/X _22425_/X _22847_/X VGND VGND VPWR VPWR _22849_/A sky130_fd_sc_hd__o22a_4
XANTENNA__23370__D HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _12600_/X VGND VGND VPWR VPWR _12602_/A sky130_fd_sc_hd__buf_2
XFILLER_77_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13581_ _13831_/A _14592_/A _13580_/Y _14570_/A VGND VGND VPWR VPWR _13581_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ _12440_/C _22489_/X _24261_/Q _21045_/X VGND VGND VPWR VPWR _22779_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ _25407_/Q VGND VGND VPWR VPWR _12609_/A sky130_fd_sc_hd__inv_2
X_15320_ _15309_/A _15331_/A _15310_/B _15308_/X VGND VGND VPWR VPWR _15320_/X sky130_fd_sc_hd__or4_4
XFILLER_13_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24518_ _24465_/CLK _16584_/X HRESETn VGND VGND VPWR VPWR _24518_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25498_ _25497_/CLK _25498_/D HRESETn VGND VGND VPWR VPWR _11916_/A sky130_fd_sc_hd__dfrtp_4
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12463_ _12430_/A _12461_/A VGND VGND VPWR VPWR _12464_/C sky130_fd_sc_hd__or2_4
X_15251_ _15262_/A _15251_/B _15251_/C _15250_/X VGND VGND VPWR VPWR _15252_/A sky130_fd_sc_hd__or4_4
X_24449_ _24462_/CLK _16760_/X HRESETn VGND VGND VPWR VPWR _15003_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16562__A _24526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14202_ _20479_/A _14199_/X _13835_/X _14201_/X VGND VGND VPWR VPWR _25196_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12556__A2 _12555_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15182_ _15166_/B _15172_/X _15174_/X _15179_/B VGND VGND VPWR VPWR _15183_/A sky130_fd_sc_hd__a211o_4
X_12394_ _12410_/A VGND VGND VPWR VPWR _12394_/X sky130_fd_sc_hd__buf_2
X_14133_ _25210_/Q _14117_/X _14119_/A _14118_/Y VGND VGND VPWR VPWR _14133_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17808__D _17751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19990_ _23535_/Q VGND VGND VPWR VPWR _19990_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14064_ _14063_/X VGND VGND VPWR VPWR _14081_/A sky130_fd_sc_hd__buf_2
X_18941_ _18939_/Y _18937_/X _18940_/X _18937_/X VGND VGND VPWR VPWR _18941_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25112__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13015_ _13001_/C _13013_/A VGND VGND VPWR VPWR _13015_/X sky130_fd_sc_hd__or2_4
X_18872_ _23934_/Q _18871_/X VGND VGND VPWR VPWR _18873_/B sky130_fd_sc_hd__or2_4
XANTENNA__21627__B _20056_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17823_ _17758_/A _17822_/X VGND VGND VPWR VPWR _17823_/Y sky130_fd_sc_hd__nand2_4
XFILLER_95_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22528__B1 _22527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17754_ _17754_/A VGND VGND VPWR VPWR _17756_/A sky130_fd_sc_hd__inv_2
X_14966_ _14966_/A VGND VGND VPWR VPWR _15249_/A sky130_fd_sc_hd__inv_2
X_16705_ _16704_/Y _16700_/X _16525_/X _16700_/X VGND VGND VPWR VPWR _24472_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21643__A _21643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13917_ _13918_/D _13912_/X _14251_/A VGND VGND VPWR VPWR _13917_/X sky130_fd_sc_hd__a21o_4
X_17685_ _17685_/A _17685_/B _17681_/X VGND VGND VPWR VPWR _17685_/X sky130_fd_sc_hd__and3_4
X_14897_ _25011_/Q VGND VGND VPWR VPWR _15067_/D sky130_fd_sc_hd__inv_2
XFILLER_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19424_ _19423_/X VGND VGND VPWR VPWR _19431_/A sky130_fd_sc_hd__inv_2
X_16636_ _16629_/Y _16634_/X _16632_/Y _16635_/Y VGND VGND VPWR VPWR _16637_/A sky130_fd_sc_hd__a211o_4
X_13848_ _25242_/Q VGND VGND VPWR VPWR _13848_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24065__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19355_ _19354_/X VGND VGND VPWR VPWR _19355_/Y sky130_fd_sc_hd__inv_2
X_16567_ _24524_/Q VGND VGND VPWR VPWR _16567_/Y sky130_fd_sc_hd__inv_2
X_13779_ _13815_/A _14219_/A VGND VGND VPWR VPWR _13779_/X sky130_fd_sc_hd__or2_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22700__B1 _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18306_ _24199_/Q VGND VGND VPWR VPWR _21173_/A sky130_fd_sc_hd__inv_2
X_15518_ _15515_/Y _15511_/X HADDR[12] _15517_/X VGND VGND VPWR VPWR _15518_/X sky130_fd_sc_hd__a2bb2o_4
X_19286_ _19683_/A _18331_/X _19219_/X VGND VGND VPWR VPWR _19287_/A sky130_fd_sc_hd__or3_4
X_16498_ _16466_/A VGND VGND VPWR VPWR _16504_/A sky130_fd_sc_hd__buf_2
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17183__B2 _17254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18237_ _18237_/A VGND VGND VPWR VPWR _18237_/X sky130_fd_sc_hd__buf_2
X_15449_ _15449_/A VGND VGND VPWR VPWR _15449_/X sky130_fd_sc_hd__buf_2
XFILLER_50_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20794__A1_N _20770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18168_ _18168_/A _20226_/A VGND VGND VPWR VPWR _18169_/C sky130_fd_sc_hd__or2_4
XANTENNA__14902__A1_N _25005_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11755__B1 _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17119_ _17050_/A _17045_/X VGND VGND VPWR VPWR _17119_/X sky130_fd_sc_hd__or2_4
X_18099_ _17963_/X _18098_/X _24233_/Q _18021_/X VGND VGND VPWR VPWR _18099_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20130_ _23483_/Q VGND VGND VPWR VPWR _22192_/B sky130_fd_sc_hd__inv_2
XFILLER_104_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22767__B1 _24858_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20061_ _20061_/A VGND VGND VPWR VPWR _20061_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16446__B1 _16366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12180__B1 _12179_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22519__B1 _22498_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24835__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23820_ _23818_/CLK _19177_/X VGND VGND VPWR VPWR _19173_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16470__A1_N _16469_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23192__B1 _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23751_ _23446_/CLK _23751_/D VGND VGND VPWR VPWR _18132_/B sky130_fd_sc_hd__dfxtp_4
X_20963_ _12143_/A _20965_/B VGND VGND VPWR VPWR _20963_/X sky130_fd_sc_hd__and2_4
XFILLER_22_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21742__B2 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22702_ _22702_/A _21220_/A VGND VGND VPWR VPWR _22702_/X sky130_fd_sc_hd__or2_4
XANTENNA__15551__A _15642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17410__A2 _17401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23682_ _23682_/CLK _23682_/D VGND VGND VPWR VPWR _23682_/Q sky130_fd_sc_hd__dfxtp_4
X_20894_ _24046_/Q _20889_/X _20893_/X VGND VGND VPWR VPWR _20894_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22087__C _22086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25421_ _25449_/CLK _25421_/D HRESETn VGND VGND VPWR VPWR _12280_/A sky130_fd_sc_hd__dfrtp_4
X_22633_ _15607_/Y _22747_/B VGND VGND VPWR VPWR _22633_/X sky130_fd_sc_hd__and2_4
XFILLER_80_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25352_ _23370_/CLK _13011_/Y HRESETn VGND VGND VPWR VPWR _12374_/A sky130_fd_sc_hd__dfrtp_4
X_22564_ _22564_/A VGND VGND VPWR VPWR _22564_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_172_0_HCLK clkbuf_7_86_0_HCLK/X VGND VGND VPWR VPWR _23545_/CLK sky130_fd_sc_hd__clkbuf_1
X_21515_ _21512_/X _21513_/X _21514_/X _25509_/Q _21428_/X VGND VGND VPWR VPWR _21516_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24303_ _25526_/CLK _17615_/X HRESETn VGND VGND VPWR VPWR _17562_/A sky130_fd_sc_hd__dfrtp_4
X_25283_ _24252_/CLK _13697_/X HRESETn VGND VGND VPWR VPWR _13676_/A sky130_fd_sc_hd__dfrtp_4
X_22495_ _16515_/Y _22493_/B VGND VGND VPWR VPWR _22495_/X sky130_fd_sc_hd__and2_4
XFILLER_103_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_29_0_HCLK clkbuf_8_29_0_HCLK/A VGND VGND VPWR VPWR _25122_/CLK sky130_fd_sc_hd__clkbuf_1
X_24234_ _23826_/CLK _24234_/D HRESETn VGND VGND VPWR VPWR _24234_/Q sky130_fd_sc_hd__dfrtp_4
X_21446_ _17706_/A VGND VGND VPWR VPWR _21452_/A sky130_fd_sc_hd__buf_2
XFILLER_119_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24165_ _24159_/CLK _18530_/Y HRESETn VGND VGND VPWR VPWR _24165_/Q sky130_fd_sc_hd__dfrtp_4
X_21377_ _21377_/A _21377_/B _21376_/X VGND VGND VPWR VPWR _21377_/X sky130_fd_sc_hd__and3_4
XANTENNA__12415__A _12244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23116_ _17239_/A _22908_/X _12749_/A _22909_/X VGND VGND VPWR VPWR _23116_/X sky130_fd_sc_hd__a2bb2o_4
X_20328_ _21968_/A _20327_/X _15766_/X _20327_/X VGND VGND VPWR VPWR _20328_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24096_ _24097_/CLK _20961_/X HRESETn VGND VGND VPWR VPWR _24096_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13499__B1 _11825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23047_ _23114_/A _23033_/X _23038_/X _23046_/X VGND VGND VPWR VPWR _23047_/X sky130_fd_sc_hd__or4_4
X_20259_ _20266_/A VGND VGND VPWR VPWR _20259_/X sky130_fd_sc_hd__buf_2
XFILLER_89_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16988__A1 _16029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24576__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14820_ _14820_/A _14819_/X VGND VGND VPWR VPWR _14820_/Y sky130_fd_sc_hd__nor2_4
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24998_ _24998_/CLK _15280_/X HRESETn VGND VGND VPWR VPWR _14975_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_91_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24505__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21463__A _21658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14751_ _14749_/X _14750_/X _14746_/X VGND VGND VPWR VPWR _25050_/D sky130_fd_sc_hd__o21a_4
XFILLER_63_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11963_ _11957_/Y _17445_/B VGND VGND VPWR VPWR _11963_/X sky130_fd_sc_hd__or2_4
X_23949_ _25098_/CLK _23949_/D HRESETn VGND VGND VPWR VPWR _20531_/A sky130_fd_sc_hd__dfstp_4
X_13702_ _13702_/A _13702_/B VGND VGND VPWR VPWR _13702_/Y sky130_fd_sc_hd__nand2_4
X_17470_ _13191_/A _17469_/X _13191_/A _17469_/X VGND VGND VPWR VPWR _17489_/B sky130_fd_sc_hd__a2bb2o_4
X_11894_ _11924_/A _11894_/B VGND VGND VPWR VPWR _11894_/X sky130_fd_sc_hd__and2_4
X_14682_ _21247_/A _14682_/B VGND VGND VPWR VPWR _14750_/A sky130_fd_sc_hd__and2_4
XFILLER_45_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16421_ _16421_/A VGND VGND VPWR VPWR _16421_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13633_ _13634_/A _13633_/B _13627_/X _13633_/D VGND VGND VPWR VPWR _13633_/X sky130_fd_sc_hd__or4_4
X_19140_ _19139_/Y _19137_/X _19071_/X _19137_/X VGND VGND VPWR VPWR _23833_/D sky130_fd_sc_hd__a2bb2o_4
X_16352_ _16352_/A VGND VGND VPWR VPWR _16352_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13564_ _13564_/A _13558_/X _13564_/C _13564_/D VGND VGND VPWR VPWR _13588_/B sky130_fd_sc_hd__or4_4
XFILLER_73_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15303_ _15390_/A _15389_/A _15388_/C _15092_/Y VGND VGND VPWR VPWR _15303_/X sky130_fd_sc_hd__or4_4
X_12515_ _25415_/Q VGND VGND VPWR VPWR _12645_/A sky130_fd_sc_hd__inv_2
X_19071_ _16781_/X VGND VGND VPWR VPWR _19071_/X sky130_fd_sc_hd__buf_2
X_13495_ _16183_/A _13468_/X VGND VGND VPWR VPWR _13495_/X sky130_fd_sc_hd__or2_4
X_16283_ _16278_/Y _16282_/X _11743_/X _16282_/X VGND VGND VPWR VPWR _24630_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25364__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18022_ _17963_/X _18020_/X _24235_/Q _18021_/X VGND VGND VPWR VPWR _24235_/D sky130_fd_sc_hd__o22a_4
XFILLER_117_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12446_ _12429_/X _12440_/X _12446_/C VGND VGND VPWR VPWR _12446_/X sky130_fd_sc_hd__and3_4
X_15234_ _14961_/X _15232_/A VGND VGND VPWR VPWR _15234_/X sky130_fd_sc_hd__or2_4
XFILLER_138_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12377_ _12377_/A VGND VGND VPWR VPWR _12377_/Y sky130_fd_sc_hd__inv_2
X_15165_ _15165_/A _15165_/B VGND VGND VPWR VPWR _15165_/X sky130_fd_sc_hd__or2_4
XANTENNA__19862__B1 _19797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14116_ _14116_/A _14116_/B _14102_/A VGND VGND VPWR VPWR _14117_/B sky130_fd_sc_hd__or3_4
X_15096_ _15096_/A VGND VGND VPWR VPWR _15096_/Y sky130_fd_sc_hd__inv_2
X_19973_ _19973_/A VGND VGND VPWR VPWR _19991_/A sky130_fd_sc_hd__inv_2
XFILLER_99_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18924_ _18923_/X VGND VGND VPWR VPWR _18937_/A sky130_fd_sc_hd__inv_2
XFILLER_84_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15636__A _21280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14047_ _13999_/X VGND VGND VPWR VPWR _14047_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18012__A _18184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16428__B1 _16340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18855_ _24540_/Q _18782_/X _16510_/Y _18789_/A VGND VGND VPWR VPWR _18855_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16979__A1 _24710_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16979__B2 _17038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17806_ _17806_/A VGND VGND VPWR VPWR _24267_/D sky130_fd_sc_hd__inv_2
XFILLER_67_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18786_ _18623_/Y _18782_/X _18786_/C _18786_/D VGND VGND VPWR VPWR _18792_/C sky130_fd_sc_hd__or4_4
X_15998_ _15990_/Y _15997_/X _11743_/X _15997_/X VGND VGND VPWR VPWR _24734_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23174__B1 _22997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24246__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17737_ _16953_/X VGND VGND VPWR VPWR _17737_/X sky130_fd_sc_hd__buf_2
X_14949_ _25009_/Q VGND VGND VPWR VPWR _14949_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_5_20_0_HCLK_A clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12465__A1 _12235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17668_ _17517_/Y _17674_/B VGND VGND VPWR VPWR _17672_/B sky130_fd_sc_hd__or2_4
XFILLER_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19407_ _18996_/X VGND VGND VPWR VPWR _19407_/X sky130_fd_sc_hd__buf_2
XFILLER_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16619_ _16618_/Y _16614_/X _16442_/X _16614_/X VGND VGND VPWR VPWR _24504_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17599_ _17611_/A _17837_/A VGND VGND VPWR VPWR _17600_/D sky130_fd_sc_hd__and2_4
XFILLER_50_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19338_ _18045_/B VGND VGND VPWR VPWR _19338_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_245_0_HCLK clkbuf_8_245_0_HCLK/A VGND VGND VPWR VPWR _25016_/CLK sky130_fd_sc_hd__clkbuf_1
X_19269_ _22205_/B _19266_/X _16867_/X _19266_/X VGND VGND VPWR VPWR _19269_/X sky130_fd_sc_hd__a2bb2o_4
X_21300_ _21280_/B _21294_/X _21296_/X _24704_/Q _21299_/X VGND VGND VPWR VPWR _21300_/X
+ sky130_fd_sc_hd__a32o_4
X_22280_ _22280_/A VGND VGND VPWR VPWR _22280_/X sky130_fd_sc_hd__buf_2
XFILLER_117_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25034__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21231_ _21253_/A _21231_/B VGND VGND VPWR VPWR _21231_/X sky130_fd_sc_hd__or2_4
XANTENNA__19853__B1 _19783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16667__B1 _16398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21162_ _21162_/A VGND VGND VPWR VPWR _21162_/X sky130_fd_sc_hd__buf_2
XANTENNA__21660__B1 _18299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20113_ _23489_/Q VGND VGND VPWR VPWR _21892_/B sky130_fd_sc_hd__inv_2
XANTENNA__12566__A2_N _24854_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15546__A _22915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21093_ _21040_/A _21086_/X _21093_/C VGND VGND VPWR VPWR _21093_/X sky130_fd_sc_hd__and3_4
XFILLER_132_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19605__B1 _19462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20044_ _20044_/A VGND VGND VPWR VPWR _20057_/A sky130_fd_sc_hd__inv_2
XFILLER_131_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24921_ _23550_/CLK _24921_/D HRESETn VGND VGND VPWR VPWR _15523_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_28_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24852_ _24852_/CLK _15755_/X HRESETn VGND VGND VPWR VPWR _24852_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23803_ _23798_/CLK _19225_/X VGND VGND VPWR VPWR _13211_/B sky130_fd_sc_hd__dfxtp_4
X_21995_ _21995_/A VGND VGND VPWR VPWR _21995_/Y sky130_fd_sc_hd__inv_2
X_24783_ _24821_/CLK _24783_/D HRESETn VGND VGND VPWR VPWR _24783_/Q sky130_fd_sc_hd__dfrtp_4
X_20946_ _13667_/C VGND VGND VPWR VPWR _20946_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23734_ _23722_/CLK _23734_/D VGND VGND VPWR VPWR _18171_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_121_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23969__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _20879_/A VGND VGND VPWR VPWR _20877_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12208__B2 _12207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_55_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23665_ _24930_/CLK _23665_/D VGND VGND VPWR VPWR _19621_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25404_ _25400_/CLK _25404_/D HRESETn VGND VGND VPWR VPWR _12520_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22616_ _17249_/Y _22534_/X _22615_/Y VGND VGND VPWR VPWR _22616_/X sky130_fd_sc_hd__o21a_4
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23596_ _23434_/CLK _23596_/D VGND VGND VPWR VPWR _19821_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22140__A1 _24708_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22547_ _21066_/A VGND VGND VPWR VPWR _22547_/X sky130_fd_sc_hd__buf_2
X_25335_ _25351_/CLK _13076_/X HRESETn VGND VGND VPWR VPWR _25335_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22691__A2 _21587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12300_ _12299_/Y _24832_/Q _12299_/Y _24832_/Q VGND VGND VPWR VPWR _12300_/X sky130_fd_sc_hd__a2bb2o_4
X_13280_ _13386_/A _13280_/B _13280_/C VGND VGND VPWR VPWR _13285_/B sky130_fd_sc_hd__and3_4
X_22478_ _22478_/A _22626_/B VGND VGND VPWR VPWR _22478_/X sky130_fd_sc_hd__or2_4
X_25266_ _25055_/CLK _13764_/X HRESETn VGND VGND VPWR VPWR _13754_/A sky130_fd_sc_hd__dfrtp_4
X_12231_ _21433_/A VGND VGND VPWR VPWR _12231_/Y sky130_fd_sc_hd__inv_2
X_21429_ _16640_/A _21426_/X _21427_/X _11860_/A _21428_/X VGND VGND VPWR VPWR _21429_/X
+ sky130_fd_sc_hd__a32o_4
X_24217_ _25279_/CLK _24217_/D HRESETn VGND VGND VPWR VPWR _21967_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22443__A2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25197_ _25098_/CLK _14184_/Y HRESETn VGND VGND VPWR VPWR _25197_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12162_ _12157_/X VGND VGND VPWR VPWR _12163_/B sky130_fd_sc_hd__inv_2
XANTENNA__21458__A _21458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16992__A1_N _24720_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24148_ _24148_/CLK _24148_/D HRESETn VGND VGND VPWR VPWR _24148_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24757__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12093_ _13789_/B VGND VGND VPWR VPWR _12093_/X sky130_fd_sc_hd__buf_2
X_16970_ _16075_/Y _17043_/A _16075_/Y _17043_/A VGND VGND VPWR VPWR _16971_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24079_ _23995_/CLK _24079_/D HRESETn VGND VGND VPWR VPWR _20443_/A sky130_fd_sc_hd__dfrtp_4
X_15921_ _15677_/X _15920_/Y _15684_/A _15920_/Y VGND VGND VPWR VPWR _15921_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22746__A3 _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18640_ _18809_/A VGND VGND VPWR VPWR _18680_/B sky130_fd_sc_hd__inv_2
XFILLER_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15852_ _15852_/A VGND VGND VPWR VPWR _15852_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14803_ _14817_/C _14803_/B _14803_/C VGND VGND VPWR VPWR _14804_/A sky130_fd_sc_hd__or3_4
X_18571_ _18416_/Y _18574_/B VGND VGND VPWR VPWR _18571_/Y sky130_fd_sc_hd__nand2_4
X_15783_ _15782_/X VGND VGND VPWR VPWR _15784_/B sky130_fd_sc_hd__buf_2
X_12995_ _12995_/A _12363_/Y _13106_/A _12311_/Y VGND VGND VPWR VPWR _12995_/X sky130_fd_sc_hd__or4_4
XANTENNA__22903__B1 _25526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17522_ _25525_/Q _24296_/Q _11787_/Y _17521_/Y VGND VGND VPWR VPWR _17522_/X sky130_fd_sc_hd__o22a_4
X_14734_ _25055_/Q VGND VGND VPWR VPWR _14734_/Y sky130_fd_sc_hd__inv_2
X_11946_ _19629_/A VGND VGND VPWR VPWR _11946_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17453_ _17453_/A _17453_/B VGND VGND VPWR VPWR _17456_/A sky130_fd_sc_hd__and2_4
X_14665_ _18972_/A VGND VGND VPWR VPWR _14665_/X sky130_fd_sc_hd__buf_2
XFILLER_44_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11877_ _11877_/A _11876_/X VGND VGND VPWR VPWR _11878_/B sky130_fd_sc_hd__and2_4
X_16404_ _15147_/Y _16400_/X _16403_/X _16400_/X VGND VGND VPWR VPWR _24587_/D sky130_fd_sc_hd__a2bb2o_4
X_13616_ _17995_/A VGND VGND VPWR VPWR _18057_/A sky130_fd_sc_hd__buf_2
X_17384_ _17242_/A _17384_/B VGND VGND VPWR VPWR _17384_/X sky130_fd_sc_hd__or2_4
X_14596_ _14559_/Y _14596_/B VGND VGND VPWR VPWR _14596_/Y sky130_fd_sc_hd__nand2_4
X_19123_ _19122_/Y _19120_/X _19056_/X _19120_/X VGND VGND VPWR VPWR _19123_/X sky130_fd_sc_hd__a2bb2o_4
X_16335_ _16334_/Y _16330_/X _16238_/X _16330_/X VGND VGND VPWR VPWR _16335_/X sky130_fd_sc_hd__a2bb2o_4
X_13547_ _22612_/A _14558_/A _22612_/A _14558_/A VGND VGND VPWR VPWR _13554_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22682__A2 _23126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18007__A _18087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19054_ _23862_/Q VGND VGND VPWR VPWR _19054_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16453__C _15533_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16266_ _14470_/A VGND VGND VPWR VPWR _16266_/X sky130_fd_sc_hd__buf_2
X_13478_ _13474_/Y _13477_/X _11833_/X _13477_/X VGND VGND VPWR VPWR _25311_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_12_0_HCLK clkbuf_7_6_0_HCLK/X VGND VGND VPWR VPWR _23496_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18005_ _18005_/A _18002_/X _18005_/C VGND VGND VPWR VPWR _18006_/C sky130_fd_sc_hd__and3_4
X_15217_ _15212_/A _15211_/X _15199_/X _15214_/B VGND VGND VPWR VPWR _15218_/A sky130_fd_sc_hd__a211o_4
XFILLER_86_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12429_ _12509_/A VGND VGND VPWR VPWR _12429_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_75_0_HCLK clkbuf_8_75_0_HCLK/A VGND VGND VPWR VPWR _25178_/CLK sky130_fd_sc_hd__clkbuf_1
X_16197_ _23200_/A VGND VGND VPWR VPWR _16197_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16649__B1 _16380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12922__A2 _12903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15148_ _15087_/Y _24593_/Q _24983_/Q _15147_/Y VGND VGND VPWR VPWR _15152_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24498__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15079_ _24969_/Q _15077_/Y _15331_/A _15090_/A VGND VGND VPWR VPWR _15079_/X sky130_fd_sc_hd__a2bb2o_4
X_19956_ _23546_/Q VGND VGND VPWR VPWR _22016_/B sky130_fd_sc_hd__inv_2
XANTENNA__24427__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18907_ _18901_/Y VGND VGND VPWR VPWR _18907_/X sky130_fd_sc_hd__buf_2
XFILLER_68_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19887_ _19887_/A VGND VGND VPWR VPWR _19887_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18838_ _18838_/A _18838_/B _18836_/X _18837_/X VGND VGND VPWR VPWR _18838_/X sky130_fd_sc_hd__or4_4
XFILLER_68_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24080__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16821__B1 HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18769_ _18759_/A _18767_/X _18768_/X VGND VGND VPWR VPWR _24128_/D sky130_fd_sc_hd__and3_4
XANTENNA__12438__A1 _12433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20800_ _20799_/Y _20800_/B VGND VGND VPWR VPWR _20800_/X sky130_fd_sc_hd__and2_4
XFILLER_36_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21780_ _22531_/B _21779_/X _13572_/Y _22531_/B VGND VGND VPWR VPWR _21780_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22927__A _22927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20731_ _13133_/B VGND VGND VPWR VPWR _20731_/Y sky130_fd_sc_hd__inv_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20920__A2 _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25286__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23450_ _23660_/CLK _20218_/X VGND VGND VPWR VPWR _20216_/A sky130_fd_sc_hd__dfxtp_4
X_20662_ _20662_/A _20662_/B VGND VGND VPWR VPWR _20662_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__17535__A2_N _24295_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22122__A1 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22401_ _22265_/X _22400_/X _22130_/C _24814_/Q _22268_/X VGND VGND VPWR VPWR _22401_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_17_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11949__B1 _11948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22122__B2 _21533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23381_ _24219_/CLK _20392_/X VGND VGND VPWR VPWR _23381_/Q sky130_fd_sc_hd__dfxtp_4
X_20593_ _20447_/A _20591_/X _20592_/Y VGND VGND VPWR VPWR _20593_/X sky130_fd_sc_hd__and3_4
XFILLER_52_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15539__A1_N _13789_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22332_ _21944_/A _22332_/B VGND VGND VPWR VPWR _22332_/X sky130_fd_sc_hd__or2_4
XANTENNA__11868__A1_N _11864_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25120_ _25122_/CLK _25120_/D HRESETn VGND VGND VPWR VPWR _14446_/A sky130_fd_sc_hd__dfstp_4
X_25051_ _24089_/CLK _14747_/X HRESETn VGND VGND VPWR VPWR _21403_/A sky130_fd_sc_hd__dfrtp_4
X_22263_ _22263_/A VGND VGND VPWR VPWR _22293_/B sky130_fd_sc_hd__inv_2
XANTENNA__18629__A1 _24531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18629__B2 _18705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24002_ _24033_/CLK _20702_/Y HRESETn VGND VGND VPWR VPWR _20699_/A sky130_fd_sc_hd__dfrtp_4
X_21214_ _16719_/Y _21859_/B VGND VGND VPWR VPWR _21220_/B sky130_fd_sc_hd__or2_4
X_22194_ _22193_/X _22194_/B VGND VGND VPWR VPWR _22194_/X sky130_fd_sc_hd__or2_4
XFILLER_104_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24850__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21145_ _14241_/Y _14220_/A _17436_/Y _21355_/A VGND VGND VPWR VPWR _21145_/X sky130_fd_sc_hd__o22a_4
XFILLER_133_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21076_ _21075_/X VGND VGND VPWR VPWR _21076_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20027_ _22253_/B _20024_/X _19978_/X _20024_/X VGND VGND VPWR VPWR _23523_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11806__A1_N _11802_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24904_ _24049_/CLK _15578_/X HRESETn VGND VGND VPWR VPWR _15577_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16812__B1 HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24835_ _24832_/CLK _24835_/D HRESETn VGND VGND VPWR VPWR _12364_/A sky130_fd_sc_hd__dfrtp_4
X_11800_ _11800_/A VGND VGND VPWR VPWR _11800_/X sky130_fd_sc_hd__buf_2
X_12780_ _12778_/A _22895_/A _12850_/C _12779_/Y VGND VGND VPWR VPWR _12780_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11970__C _11970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24766_ _24766_/CLK _24766_/D HRESETn VGND VGND VPWR VPWR _24766_/Q sky130_fd_sc_hd__dfrtp_4
X_21978_ _22389_/A _21978_/B _21978_/C _23408_/Q VGND VGND VPWR VPWR _21978_/X sky130_fd_sc_hd__or4_4
XFILLER_15_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21741__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11731_ _24920_/Q _13777_/A _11731_/C _11731_/D VGND VGND VPWR VPWR _11732_/A sky130_fd_sc_hd__or4_4
XPHY_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23717_ _23722_/CLK _19465_/X VGND VGND VPWR VPWR _18206_/B sky130_fd_sc_hd__dfxtp_4
X_20929_ _20931_/A VGND VGND VPWR VPWR _20929_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24697_ _24699_/CLK _16095_/X HRESETn VGND VGND VPWR VPWR _16092_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14450_ _14177_/Y _14448_/X _14239_/X _14448_/X VGND VGND VPWR VPWR _25118_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _25274_/Q _11661_/Y _11656_/Y _21967_/A VGND VGND VPWR VPWR _11662_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23648_ _23649_/CLK _19674_/X VGND VGND VPWR VPWR _19673_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_109_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _17452_/B _13401_/B VGND VGND VPWR VPWR _13403_/B sky130_fd_sc_hd__or2_4
XANTENNA__25180__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14381_ _14381_/A _14394_/B VGND VGND VPWR VPWR _14383_/A sky130_fd_sc_hd__nor2_4
XANTENNA__20124__B1 _20123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23579_ _23388_/CLK _19871_/X VGND VGND VPWR VPWR _23579_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16120_ _22865_/A VGND VGND VPWR VPWR _16120_/Y sky130_fd_sc_hd__inv_2
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13332_ _13461_/A _13326_/X _13331_/X VGND VGND VPWR VPWR _13332_/X sky130_fd_sc_hd__or3_4
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25318_ _23377_/CLK _13296_/X HRESETn VGND VGND VPWR VPWR _25318_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16051_ _24712_/Q VGND VGND VPWR VPWR _16051_/Y sky130_fd_sc_hd__inv_2
X_13263_ _13402_/A _13263_/B VGND VGND VPWR VPWR _13263_/X sky130_fd_sc_hd__or2_4
X_25249_ _25290_/CLK _13836_/X HRESETn VGND VGND VPWR VPWR _13557_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15002_ _15002_/A _15002_/B _14999_/X _15002_/D VGND VGND VPWR VPWR _15002_/X sky130_fd_sc_hd__or4_4
X_12214_ _22892_/A VGND VGND VPWR VPWR _12214_/Y sky130_fd_sc_hd__inv_2
X_13194_ _11963_/X _11974_/X VGND VGND VPWR VPWR _13194_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24591__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12145_ _12135_/X _12136_/X _12140_/X _12145_/D VGND VGND VPWR VPWR _12145_/X sky130_fd_sc_hd__or4_4
X_19810_ _13330_/B VGND VGND VPWR VPWR _19810_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15186__A _25022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12117__B1 _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24520__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12076_ _12076_/A VGND VGND VPWR VPWR _12076_/Y sky130_fd_sc_hd__inv_2
X_16953_ _16953_/A _16952_/X VGND VGND VPWR VPWR _16953_/X sky130_fd_sc_hd__or2_4
X_19741_ _19739_/Y _19735_/X _19740_/X _19735_/X VGND VGND VPWR VPWR _19741_/X sky130_fd_sc_hd__a2bb2o_4
X_15904_ _15900_/A VGND VGND VPWR VPWR _15904_/X sky130_fd_sc_hd__buf_2
X_19672_ _19671_/Y _19669_/X _19547_/X _19669_/X VGND VGND VPWR VPWR _23649_/D sky130_fd_sc_hd__a2bb2o_4
X_16884_ _19797_/A VGND VGND VPWR VPWR _16884_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18623_ _18623_/A VGND VGND VPWR VPWR _18623_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16803__B1 HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15835_ _15819_/A VGND VGND VPWR VPWR _15835_/X sky130_fd_sc_hd__buf_2
XANTENNA__13434__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18554_ _18467_/Y _18552_/A VGND VGND VPWR VPWR _18554_/X sky130_fd_sc_hd__or2_4
X_15766_ _15766_/A VGND VGND VPWR VPWR _15766_/X sky130_fd_sc_hd__buf_2
X_12978_ _25355_/Q _12631_/B VGND VGND VPWR VPWR _12978_/X sky130_fd_sc_hd__or2_4
XFILLER_75_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17505_ _17505_/A _17505_/B _17505_/C _17504_/X VGND VGND VPWR VPWR _17505_/X sky130_fd_sc_hd__or4_4
XFILLER_33_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14717_ _13735_/A _13759_/A _25267_/Q _13759_/Y VGND VGND VPWR VPWR _14717_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18020__A2 _17994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11929_ _19615_/A VGND VGND VPWR VPWR _11929_/Y sky130_fd_sc_hd__inv_2
X_18485_ _18517_/A _18485_/B _18484_/Y VGND VGND VPWR VPWR _18485_/X sky130_fd_sc_hd__and3_4
X_15697_ _15680_/A _15691_/Y _15687_/C _15696_/X VGND VGND VPWR VPWR _15697_/X sky130_fd_sc_hd__o22a_4
XFILLER_127_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17436_ _17436_/A VGND VGND VPWR VPWR _17436_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14648_ _18005_/A VGND VGND VPWR VPWR _14648_/X sky130_fd_sc_hd__buf_2
XFILLER_60_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22104__A1 _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17367_ _17349_/A _17370_/B _17271_/X VGND VGND VPWR VPWR _17367_/Y sky130_fd_sc_hd__a21oi_4
X_14579_ _14558_/X _14579_/B VGND VGND VPWR VPWR _14582_/B sky130_fd_sc_hd__and2_4
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19106_ _19106_/A VGND VGND VPWR VPWR _19106_/Y sky130_fd_sc_hd__inv_2
X_16318_ _22860_/A VGND VGND VPWR VPWR _16318_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17298_ _17293_/A _17293_/B _17279_/X _17295_/B VGND VGND VPWR VPWR _17298_/X sky130_fd_sc_hd__a211o_4
X_19037_ _19152_/D VGND VGND VPWR VPWR _19038_/B sky130_fd_sc_hd__buf_2
XFILLER_51_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16899__A1_N _22556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24679__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16249_ _16249_/A VGND VGND VPWR VPWR _16249_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24608__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16822__A1_N _14941_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12108__B1 _11833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24261__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19939_ _19938_/Y _19936_/X _19622_/X _19936_/X VGND VGND VPWR VPWR _19939_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15824__A _22873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22950_ _24453_/Q _23019_/B _23019_/C VGND VGND VPWR VPWR _22950_/X sky130_fd_sc_hd__and3_4
XANTENNA__22591__A1 _22476_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22591__B2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21901_ _21601_/A _21901_/B _21901_/C VGND VGND VPWR VPWR _21901_/X sky130_fd_sc_hd__and3_4
XFILLER_3_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22881_ _24520_/Q _21067_/A _22797_/X _22880_/X VGND VGND VPWR VPWR _22882_/C sky130_fd_sc_hd__a211o_4
XANTENNA__25467__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12886__C _12600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_120_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_241_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24620_ _24346_/CLK _24620_/D HRESETn VGND VGND VPWR VPWR _22971_/A sky130_fd_sc_hd__dfrtp_4
X_21832_ _14207_/Y _14195_/B _14266_/Y _14258_/A VGND VGND VPWR VPWR _21832_/X sky130_fd_sc_hd__o22a_4
XFILLER_83_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11792__A1_N _11790_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21561__A _12096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21763_ _21763_/A _21763_/B _21762_/X VGND VGND VPWR VPWR _21763_/X sky130_fd_sc_hd__and3_4
X_24551_ _24553_/CLK _16496_/X HRESETn VGND VGND VPWR VPWR _24551_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20714_ _20712_/A _20707_/X _20713_/X VGND VGND VPWR VPWR _20714_/Y sky130_fd_sc_hd__a21oi_4
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23502_ _24208_/CLK _23502_/D VGND VGND VPWR VPWR _13412_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21280__B _21280_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21694_ _24775_/Q _22998_/A VGND VGND VPWR VPWR _21694_/X sky130_fd_sc_hd__or2_4
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24482_ _24413_/CLK _16681_/X HRESETn VGND VGND VPWR VPWR _24482_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15478__A1_N _14868_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11799__A HWDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20645_ _20645_/A VGND VGND VPWR VPWR _23977_/D sky130_fd_sc_hd__inv_2
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23433_ _23609_/CLK _23433_/D VGND VGND VPWR VPWR _23433_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23364_ _21007_/X VGND VGND VPWR VPWR IRQ[10] sky130_fd_sc_hd__buf_2
X_20576_ _14423_/Y _20556_/X _20546_/X _20575_/X VGND VGND VPWR VPWR _20577_/A sky130_fd_sc_hd__a211o_4
XFILLER_20_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17522__A1 _25525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25103_ _25178_/CLK _25103_/D HRESETn VGND VGND VPWR VPWR _25103_/Q sky130_fd_sc_hd__dfrtp_4
X_22315_ _22314_/X VGND VGND VPWR VPWR _22315_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23295_ _16378_/A _23327_/B VGND VGND VPWR VPWR _23295_/X sky130_fd_sc_hd__or2_4
XFILLER_69_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24349__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22246_ _22246_/A _22246_/B VGND VGND VPWR VPWR _22246_/X sky130_fd_sc_hd__or2_4
XANTENNA__21606__B1 _14712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25034_ _25029_/CLK _14857_/X HRESETn VGND VGND VPWR VPWR _14814_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_106_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21082__A1 _24807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22177_ _20500_/A _21843_/X _23962_/Q _21351_/B VGND VGND VPWR VPWR _22177_/X sky130_fd_sc_hd__a2bb2o_4
X_21128_ _25452_/Q _12093_/X _12046_/Y _12093_/X VGND VGND VPWR VPWR _21128_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13847__B1 _13515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13950_ _13970_/A _13944_/Y _13950_/C _13949_/X VGND VGND VPWR VPWR _13950_/X sky130_fd_sc_hd__or4_4
X_21059_ _21040_/A _21059_/B _21059_/C VGND VGND VPWR VPWR _21059_/X sky130_fd_sc_hd__and3_4
XFILLER_47_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19206__A _16781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12901_ _12979_/A VGND VGND VPWR VPWR _12936_/A sky130_fd_sc_hd__buf_2
XFILLER_19_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23984__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13881_ _13871_/X _13880_/X _14273_/A _13856_/Y VGND VGND VPWR VPWR _25232_/D sky130_fd_sc_hd__o22a_4
XFILLER_46_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15620_ _16057_/A VGND VGND VPWR VPWR _15620_/X sky130_fd_sc_hd__buf_2
X_12832_ _25383_/Q _12820_/Y _12819_/X _24776_/Q VGND VGND VPWR VPWR _12832_/X sky130_fd_sc_hd__a2bb2o_4
X_24818_ _24842_/CLK _24818_/D HRESETn VGND VGND VPWR VPWR _24818_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14272__B1 _13803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25137__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15551_ _15642_/A _15551_/B VGND VGND VPWR VPWR _15777_/A sky130_fd_sc_hd__or2_4
XFILLER_15_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12763_ _12754_/X _12757_/X _12760_/X _12763_/D VGND VGND VPWR VPWR _12763_/X sky130_fd_sc_hd__or4_4
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24749_ _24785_/CLK _24749_/D HRESETn VGND VGND VPWR VPWR _24749_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _23951_/Q VGND VGND VPWR VPWR _14502_/X sky130_fd_sc_hd__buf_2
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _24061_/Q VGND VGND VPWR VPWR _11714_/Y sky130_fd_sc_hd__inv_2
X_18270_ _13780_/X VGND VGND VPWR VPWR _18270_/X sky130_fd_sc_hd__buf_2
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _24937_/Q _15438_/X _15435_/X VGND VGND VPWR VPWR _24937_/D sky130_fd_sc_hd__a21bo_4
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12565_/Y _12693_/X VGND VGND VPWR VPWR _12695_/A sky130_fd_sc_hd__or2_4
XFILLER_15_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_25_0_HCLK clkbuf_4_12_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _16295_/Y _17236_/A _22940_/A _17220_/Y VGND VGND VPWR VPWR _17221_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14433_/A VGND VGND VPWR VPWR _21352_/A sky130_fd_sc_hd__buf_2
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15772__B1 _24842_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17152_ _17044_/B _17128_/X _17149_/Y _17067_/X VGND VGND VPWR VPWR _17153_/A sky130_fd_sc_hd__a211o_4
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14364_ _25145_/Q _14351_/X _25144_/Q _14356_/X VGND VGND VPWR VPWR _14364_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17513__A1 _11831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20815__A _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16103_ _24693_/Q VGND VGND VPWR VPWR _16103_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24772__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13315_ _13297_/X _13306_/X _13315_/C VGND VGND VPWR VPWR _13315_/X sky130_fd_sc_hd__and3_4
XANTENNA__16621__A2_N _16545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17083_ _17064_/A _17079_/X _17082_/Y VGND VGND VPWR VPWR _17083_/X sky130_fd_sc_hd__and3_4
XFILLER_6_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14295_ _14299_/A VGND VGND VPWR VPWR _14296_/B sky130_fd_sc_hd__buf_2
XFILLER_100_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24701__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16034_ _15995_/X VGND VGND VPWR VPWR _16060_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13246_ _13234_/A VGND VGND VPWR VPWR _13246_/X sky130_fd_sc_hd__buf_2
XFILLER_124_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24019__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13177_ _13177_/A VGND VGND VPWR VPWR _13177_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_149_0_HCLK clkbuf_7_74_0_HCLK/X VGND VGND VPWR VPWR _24346_/CLK sky130_fd_sc_hd__clkbuf_1
X_12128_ _12128_/A _12128_/B VGND VGND VPWR VPWR _12147_/B sky130_fd_sc_hd__and2_4
XFILLER_112_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17985_ _18168_/A _17985_/B VGND VGND VPWR VPWR _17986_/C sky130_fd_sc_hd__or2_4
XANTENNA__13838__B1 _13837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12059_ _15662_/B VGND VGND VPWR VPWR _12059_/X sky130_fd_sc_hd__buf_2
X_16936_ _16128_/Y _17754_/A _16128_/Y _17754_/A VGND VGND VPWR VPWR _16936_/X sky130_fd_sc_hd__a2bb2o_4
X_19724_ _19723_/Y _19720_/X _19700_/X _19720_/X VGND VGND VPWR VPWR _23630_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19563__A2_N _19562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22573__A1 _24412_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16867_ _19780_/A VGND VGND VPWR VPWR _16867_/X sky130_fd_sc_hd__buf_2
X_19655_ _23654_/Q VGND VGND VPWR VPWR _19655_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18955__A _16781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15818_ _15816_/X _15795_/X _15739_/X _24823_/Q _15817_/X VGND VGND VPWR VPWR _15818_/X
+ sky130_fd_sc_hd__a32o_4
X_18606_ _16581_/Y _24129_/Q _16581_/Y _24129_/Q VGND VGND VPWR VPWR _18616_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19586_ _13771_/X _24065_/Q _13775_/X _19586_/D VGND VGND VPWR VPWR _19587_/A sky130_fd_sc_hd__and4_4
X_16798_ _16794_/Y _16797_/X _16376_/X _16797_/X VGND VGND VPWR VPWR _16798_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18537_ _18540_/A _18540_/B VGND VGND VPWR VPWR _18541_/B sky130_fd_sc_hd__or2_4
XFILLER_80_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15749_ _15728_/A VGND VGND VPWR VPWR _15749_/X sky130_fd_sc_hd__buf_2
XANTENNA__20336__B1 _19771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22876__A2 _21106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18468_ _24157_/Q VGND VGND VPWR VPWR _18468_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20887__B2 _20886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17419_ _20662_/A _17417_/X _17418_/X _17417_/X VGND VGND VPWR VPWR _17419_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19501__A2_N _19495_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18399_ _22539_/A _18566_/A _16199_/Y _24171_/Q VGND VGND VPWR VPWR _18399_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_14_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12508__A _21065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20430_ _20426_/B VGND VGND VPWR VPWR _20447_/A sky130_fd_sc_hd__buf_2
XFILLER_105_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13834__A1_N _13575_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22643__C _22622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20361_ _20360_/Y VGND VGND VPWR VPWR _20361_/X sky130_fd_sc_hd__buf_2
XFILLER_119_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22100_ _14480_/Y _21548_/B _25094_/Q _22111_/B VGND VGND VPWR VPWR _22101_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24442__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23080_ _21409_/A _23078_/Y _22826_/X _23079_/X VGND VGND VPWR VPWR _23081_/A sky130_fd_sc_hd__o22a_4
X_20292_ _23421_/Q VGND VGND VPWR VPWR _20292_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_45_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22031_ _22025_/A _22027_/X _22028_/X _22029_/X _22030_/X VGND VGND VPWR VPWR _22031_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_88_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22800__A2 _21067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21556__A _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23982_ _24942_/CLK _20662_/Y HRESETn VGND VGND VPWR VPWR _23982_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22933_ _23002_/A _22920_/Y _22926_/X _22933_/D VGND VGND VPWR VPWR _22933_/X sky130_fd_sc_hd__or4_4
XFILLER_84_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22864_ _22654_/A VGND VGND VPWR VPWR _22864_/X sky130_fd_sc_hd__buf_2
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24603_ _24600_/CLK _24603_/D HRESETn VGND VGND VPWR VPWR _21852_/A sky130_fd_sc_hd__dfrtp_4
X_21815_ _21799_/X _21814_/X _21493_/X VGND VGND VPWR VPWR _21815_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_25_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22795_ _22795_/A VGND VGND VPWR VPWR _23002_/A sky130_fd_sc_hd__buf_2
XFILLER_19_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24534_ _24502_/CLK _24534_/D HRESETn VGND VGND VPWR VPWR _24534_/Q sky130_fd_sc_hd__dfrtp_4
X_21746_ _21623_/A _19253_/Y VGND VGND VPWR VPWR _21746_/X sky130_fd_sc_hd__or2_4
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24465_ _24465_/CLK _24465_/D HRESETn VGND VGND VPWR VPWR _24465_/Q sky130_fd_sc_hd__dfrtp_4
X_21677_ _21648_/A _19627_/Y VGND VGND VPWR VPWR _21678_/C sky130_fd_sc_hd__or2_4
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12568__B1 _12567_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23416_ _23714_/CLK _23416_/D VGND VGND VPWR VPWR _23416_/Q sky130_fd_sc_hd__dfxtp_4
X_20628_ _20604_/Y VGND VGND VPWR VPWR _20628_/X sky130_fd_sc_hd__buf_2
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19496__B2 _19495_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24396_ _24396_/CLK _24396_/D HRESETn VGND VGND VPWR VPWR _20092_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23011__A _22270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20559_ _22302_/A _20556_/X _20547_/X _20558_/X VGND VGND VPWR VPWR _20560_/A sky130_fd_sc_hd__a211o_4
XANTENNA__15729__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23347_ VGND VGND VPWR VPWR _23347_/HI IRQ[13] sky130_fd_sc_hd__conb_1
X_13100_ _13084_/B _13100_/B _13115_/C VGND VGND VPWR VPWR _25328_/D sky130_fd_sc_hd__and3_4
XFILLER_138_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24183__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14080_ _23993_/Q _14069_/X _14073_/X _13990_/C _14076_/X VGND VGND VPWR VPWR _14080_/X
+ sky130_fd_sc_hd__a32o_4
X_23278_ _23278_/A _23310_/B VGND VGND VPWR VPWR _23278_/X sky130_fd_sc_hd__or2_4
XANTENNA__22850__A _22792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24112__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13031_ _13026_/A VGND VGND VPWR VPWR _13031_/X sky130_fd_sc_hd__buf_2
X_25017_ _25020_/CLK _15207_/Y HRESETn VGND VGND VPWR VPWR _25017_/Q sky130_fd_sc_hd__dfrtp_4
X_22229_ _22229_/A _22229_/B VGND VGND VPWR VPWR _22229_/X sky130_fd_sc_hd__or2_4
XFILLER_105_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21466__A _21658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25389__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_2_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17770_ _16953_/X _17837_/A VGND VGND VPWR VPWR _17771_/B sky130_fd_sc_hd__and2_4
X_14982_ _15267_/A _14890_/A _14981_/X _16850_/A VGND VGND VPWR VPWR _14982_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25318__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16279__B _15993_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16721_ _16719_/Y _16658_/A _16720_/X _16658_/A VGND VGND VPWR VPWR _16721_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22555__B2 _22554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13933_ _13926_/C VGND VGND VPWR VPWR _13957_/B sky130_fd_sc_hd__buf_2
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19440_ _18172_/B VGND VGND VPWR VPWR _19440_/Y sky130_fd_sc_hd__inv_2
X_16652_ _16650_/Y _16646_/X _16384_/X _16651_/X VGND VGND VPWR VPWR _24494_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18297__A1_N _21491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13864_ _20466_/B _13861_/X _13862_/Y _13863_/X VGND VGND VPWR VPWR _13864_/X sky130_fd_sc_hd__o22a_4
XFILLER_62_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15603_ _15602_/Y _15600_/X _11804_/X _15600_/X VGND VGND VPWR VPWR _15603_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12815_ _12807_/X _12815_/B _12815_/C _12814_/X VGND VGND VPWR VPWR _12815_/X sky130_fd_sc_hd__or4_4
X_19371_ _19368_/Y _19369_/X _19370_/X _19369_/X VGND VGND VPWR VPWR _23751_/D sky130_fd_sc_hd__a2bb2o_4
X_16583_ _16583_/A VGND VGND VPWR VPWR _16583_/X sky130_fd_sc_hd__buf_2
X_13795_ _16725_/A _16725_/B _13784_/C _13795_/D VGND VGND VPWR VPWR _13795_/X sky130_fd_sc_hd__and4_4
XFILLER_27_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16295__A _16295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19184__B1 _19071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18322_ _20231_/C VGND VGND VPWR VPWR _19105_/A sky130_fd_sc_hd__buf_2
X_15534_ _15533_/Y _15529_/X HADDR[5] _15529_/X VGND VGND VPWR VPWR _15534_/X sky130_fd_sc_hd__a2bb2o_4
X_12746_ _24778_/Q VGND VGND VPWR VPWR _12746_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18931__B1 _17424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18253_ _18237_/A VGND VGND VPWR VPWR _18253_/X sky130_fd_sc_hd__buf_2
XANTENNA__24953__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15465_ _24944_/Q VGND VGND VPWR VPWR _15465_/Y sky130_fd_sc_hd__inv_2
X_12677_ _12609_/A _12682_/B _12653_/X VGND VGND VPWR VPWR _12677_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ _22816_/A _17203_/Y _16352_/Y _24333_/Q VGND VGND VPWR VPWR _17204_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ _14416_/A VGND VGND VPWR VPWR _14416_/Y sky130_fd_sc_hd__inv_2
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18184_ _18184_/A _18182_/X _18184_/C VGND VGND VPWR VPWR _18184_/X sky130_fd_sc_hd__and3_4
X_15396_ _15073_/Y _15399_/B _15339_/X VGND VGND VPWR VPWR _15396_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_102_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17135_ _17041_/D _17135_/B VGND VGND VPWR VPWR _17135_/X sky130_fd_sc_hd__or2_4
XFILLER_129_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14347_ _14337_/Y _14345_/X _14346_/Y VGND VGND VPWR VPWR _14347_/X sky130_fd_sc_hd__o21a_4
XFILLER_15_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22491__B1 _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17066_ _17026_/Y _17066_/B _17025_/B _17065_/X VGND VGND VPWR VPWR _17066_/X sky130_fd_sc_hd__or4_4
XFILLER_13_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14278_ _14278_/A VGND VGND VPWR VPWR _14279_/A sky130_fd_sc_hd__buf_2
XANTENNA__22760__A _24751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16017_ _24726_/Q VGND VGND VPWR VPWR _16017_/Y sky130_fd_sc_hd__inv_2
X_13229_ _13450_/A _13226_/X _13229_/C VGND VGND VPWR VPWR _13230_/C sky130_fd_sc_hd__and3_4
XANTENNA__17854__A _17744_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17670__B1 _17590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17968_ _17975_/A VGND VGND VPWR VPWR _18204_/A sky130_fd_sc_hd__buf_2
XFILLER_85_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25059__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19707_ _19706_/Y VGND VGND VPWR VPWR _19707_/X sky130_fd_sc_hd__buf_2
X_16919_ _22484_/A _16918_/A _16142_/Y _16918_/Y VGND VGND VPWR VPWR _16922_/C sky130_fd_sc_hd__o22a_4
X_17899_ _17899_/A VGND VGND VPWR VPWR _17900_/B sky130_fd_sc_hd__inv_2
XANTENNA__17422__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19638_ _19638_/A VGND VGND VPWR VPWR _19638_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21823__B _21744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19569_ _23681_/Q VGND VGND VPWR VPWR _19569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15984__B1 _24739_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21600_ _21398_/A VGND VGND VPWR VPWR _21601_/A sky130_fd_sc_hd__buf_2
X_22580_ _17240_/Y _22534_/X _22579_/X VGND VGND VPWR VPWR _22580_/X sky130_fd_sc_hd__o21a_4
XFILLER_107_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20324__A3 _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24694__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21531_ _21531_/A _21530_/X VGND VGND VPWR VPWR _21531_/X sky130_fd_sc_hd__or2_4
XANTENNA__15736__B1 _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24623__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21462_ _21456_/A _21462_/B VGND VGND VPWR VPWR _21462_/X sky130_fd_sc_hd__or2_4
X_24250_ _24673_/CLK _24250_/D HRESETn VGND VGND VPWR VPWR _24250_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15751__A3 _15750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15154__A2_N _24570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20413_ _20411_/Y _20412_/X _20072_/X _20412_/X VGND VGND VPWR VPWR _23373_/D sky130_fd_sc_hd__a2bb2o_4
X_23201_ _24561_/Q _23166_/X _23130_/X VGND VGND VPWR VPWR _23201_/X sky130_fd_sc_hd__o21a_4
X_21393_ _21393_/A _20184_/Y VGND VGND VPWR VPWR _21394_/C sky130_fd_sc_hd__or2_4
X_24181_ _24373_/CLK _24181_/D HRESETn VGND VGND VPWR VPWR _18381_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14453__A _15851_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20344_ _20344_/A VGND VGND VPWR VPWR _22013_/B sky130_fd_sc_hd__inv_2
X_23132_ _16560_/A _22922_/X _22923_/X _23131_/X VGND VGND VPWR VPWR _23133_/C sky130_fd_sc_hd__a211o_4
XANTENNA__23026__A2 _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17764__A _17792_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23063_ _16745_/A _22998_/X _22885_/X VGND VGND VPWR VPWR _23063_/X sky130_fd_sc_hd__o21a_4
X_20275_ _23427_/Q VGND VGND VPWR VPWR _20275_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22014_ _22005_/X _22014_/B VGND VGND VPWR VPWR _22014_/X sky130_fd_sc_hd__or2_4
XANTENNA__21286__A _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20190__A _20189_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25482__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_132_0_HCLK clkbuf_7_66_0_HCLK/X VGND VGND VPWR VPWR _23854_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15284__A _15246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25411__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_195_0_HCLK clkbuf_7_97_0_HCLK/X VGND VGND VPWR VPWR _24606_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_69_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23965_ _23964_/CLK _20991_/X HRESETn VGND VGND VPWR VPWR _20995_/B sky130_fd_sc_hd__dfstp_4
XFILLER_57_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22916_ _15590_/Y _23052_/B VGND VGND VPWR VPWR _22916_/X sky130_fd_sc_hd__and2_4
XANTENNA__14227__B1 _13837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24694__CLK _25354_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23896_ _23905_/CLK _23896_/D VGND VGND VPWR VPWR _18957_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_83_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22847_ _16122_/Y _22513_/B _15931_/B _11790_/Y _22846_/X VGND VGND VPWR VPWR _22847_/X
+ sky130_fd_sc_hd__o32a_4
X_12600_ _12558_/X _12600_/B VGND VGND VPWR VPWR _12600_/X sky130_fd_sc_hd__or2_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ _13580_/A VGND VGND VPWR VPWR _13580_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22778_ _22778_/A _22778_/B _22778_/C _22777_/X VGND VGND VPWR VPWR _22778_/X sky130_fd_sc_hd__or4_4
XFILLER_38_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ _12531_/A _12525_/X _12528_/X _12530_/X VGND VGND VPWR VPWR _12558_/B sky130_fd_sc_hd__or4_4
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24517_ _24517_/CLK _24517_/D HRESETn VGND VGND VPWR VPWR _16585_/A sky130_fd_sc_hd__dfrtp_4
X_21729_ _21729_/A VGND VGND VPWR VPWR _22923_/A sky130_fd_sc_hd__buf_2
XANTENNA__15727__B1 _11767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25497_ _25497_/CLK _11927_/X HRESETn VGND VGND VPWR VPWR _11922_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24364__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15250_ _15250_/A _15267_/A _14942_/Y _15272_/A VGND VGND VPWR VPWR _15250_/X sky130_fd_sc_hd__or4_4
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12462_ _12462_/A _12461_/Y VGND VGND VPWR VPWR _12464_/B sky130_fd_sc_hd__or2_4
X_24448_ _24462_/CLK _16762_/X HRESETn VGND VGND VPWR VPWR _24448_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16038__A1_N _16037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14201_ _14201_/A VGND VGND VPWR VPWR _14201_/X sky130_fd_sc_hd__buf_2
XFILLER_71_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15181_ _15198_/A _15181_/B _15181_/C VGND VGND VPWR VPWR _25024_/D sky130_fd_sc_hd__and3_4
XANTENNA__22473__B1 _24851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12393_ _12390_/B VGND VGND VPWR VPWR _12410_/A sky130_fd_sc_hd__inv_2
XANTENNA__14950__B2 _24415_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24379_ _24720_/CLK _17104_/X HRESETn VGND VGND VPWR VPWR _24379_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14132_ _14132_/A VGND VGND VPWR VPWR _23949_/D sky130_fd_sc_hd__buf_2
XANTENNA__12961__B1 _12866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14063_ _20452_/B VGND VGND VPWR VPWR _14063_/X sky130_fd_sc_hd__buf_2
X_18940_ _14470_/A VGND VGND VPWR VPWR _18940_/X sky130_fd_sc_hd__buf_2
XFILLER_4_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13014_ _25351_/Q _13013_/Y VGND VGND VPWR VPWR _13014_/X sky130_fd_sc_hd__or2_4
X_18871_ _23933_/Q _20539_/A VGND VGND VPWR VPWR _18871_/X sky130_fd_sc_hd__or2_4
XFILLER_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_91_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17822_ _17758_/B _17825_/A VGND VGND VPWR VPWR _17822_/X sky130_fd_sc_hd__or2_4
XFILLER_58_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22528__A1 _15023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14965_ _15000_/A _14971_/A _25005_/Q _14900_/Y VGND VGND VPWR VPWR _14965_/X sky130_fd_sc_hd__a2bb2o_4
X_17753_ _24257_/Q VGND VGND VPWR VPWR _17753_/Y sky130_fd_sc_hd__inv_2
X_13916_ _13916_/A VGND VGND VPWR VPWR _14251_/A sky130_fd_sc_hd__inv_2
X_16704_ _24472_/Q VGND VGND VPWR VPWR _16704_/Y sky130_fd_sc_hd__inv_2
X_17684_ _24283_/Q _17683_/Y VGND VGND VPWR VPWR _17685_/B sky130_fd_sc_hd__or2_4
XANTENNA__21643__B _21816_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14896_ _14887_/X _14889_/X _14892_/X _14895_/X VGND VGND VPWR VPWR _14940_/A sky130_fd_sc_hd__or4_4
X_16635_ _16172_/B _16634_/B VGND VGND VPWR VPWR _16635_/Y sky130_fd_sc_hd__nor2_4
X_19423_ _19152_/A _14670_/X _14656_/Y _19152_/D VGND VGND VPWR VPWR _19423_/X sky130_fd_sc_hd__or4_4
X_13847_ _21368_/A _13843_/X _13515_/X _13843_/X VGND VGND VPWR VPWR _13847_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13442__A _13156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16566_ _16565_/Y _16563_/X _16306_/X _16563_/X VGND VGND VPWR VPWR _24525_/D sky130_fd_sc_hd__a2bb2o_4
X_19354_ _19038_/A _18987_/D _19013_/X VGND VGND VPWR VPWR _19354_/X sky130_fd_sc_hd__or3_4
X_13778_ _11733_/A _14406_/A VGND VGND VPWR VPWR _14219_/A sky130_fd_sc_hd__or2_4
X_15517_ _15535_/A VGND VGND VPWR VPWR _15517_/X sky130_fd_sc_hd__buf_2
X_18305_ _21467_/A _18303_/X _18304_/Y VGND VGND VPWR VPWR _18305_/X sky130_fd_sc_hd__o21a_4
XFILLER_128_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12729_ _12729_/A _12737_/A VGND VGND VPWR VPWR _12731_/B sky130_fd_sc_hd__or2_4
X_19285_ _19728_/A VGND VGND VPWR VPWR _19683_/A sky130_fd_sc_hd__buf_2
X_16497_ _24550_/Q VGND VGND VPWR VPWR _16497_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22474__B _22473_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22436__A1_N _17846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18236_ _18230_/B VGND VGND VPWR VPWR _18237_/A sky130_fd_sc_hd__inv_2
X_15448_ _14280_/X _24066_/Q _15441_/Y _13889_/C _15444_/X VGND VGND VPWR VPWR _15448_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17568__B _17525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24034__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18167_ _18066_/A _23766_/Q VGND VGND VPWR VPWR _18169_/B sky130_fd_sc_hd__or2_4
X_15379_ _15336_/A _15305_/C VGND VGND VPWR VPWR _15379_/X sky130_fd_sc_hd__or2_4
XFILLER_117_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17118_ _17020_/X VGND VGND VPWR VPWR _17143_/A sky130_fd_sc_hd__buf_2
XFILLER_128_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15800__A1_N _12328_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18098_ _15695_/X _18078_/X _18097_/X _24234_/Q _18019_/X VGND VGND VPWR VPWR _18098_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_89_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17049_ _17026_/Y _17066_/B VGND VGND VPWR VPWR _17050_/D sky130_fd_sc_hd__or2_4
XFILLER_131_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20060_ _20059_/Y _20057_/X _19797_/X _20057_/X VGND VGND VPWR VPWR _23510_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15815__A1_N _12341_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12180__B2 _24766_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14457__B1 _14414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_205_0_HCLK clkbuf_8_205_0_HCLK/A VGND VGND VPWR VPWR _24025_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21990__A2 _20331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23750_ _23446_/CLK _19373_/X VGND VGND VPWR VPWR _18164_/B sky130_fd_sc_hd__dfxtp_4
X_20962_ _12138_/X _12159_/X VGND VGND VPWR VPWR _24097_/D sky130_fd_sc_hd__and2_4
XFILLER_66_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24875__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22701_ _22701_/A _22698_/X _22701_/C VGND VGND VPWR VPWR _22711_/B sky130_fd_sc_hd__and3_4
XANTENNA__15551__B _15551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23681_ _24926_/CLK _19570_/X VGND VGND VPWR VPWR _23681_/Q sky130_fd_sc_hd__dfxtp_4
X_20893_ _20888_/Y _20884_/Y _20892_/Y VGND VGND VPWR VPWR _20893_/X sky130_fd_sc_hd__and3_4
XANTENNA__24804__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25420_ _25368_/CLK _12509_/X HRESETn VGND VGND VPWR VPWR _21065_/A sky130_fd_sc_hd__dfrtp_4
X_22632_ _22544_/X _22631_/X _22125_/X _25519_/Q _22922_/A VGND VGND VPWR VPWR _22632_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13432__B2 _13195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15972__A3 _11809_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25351_ _25351_/CLK _25351_/D HRESETn VGND VGND VPWR VPWR _25351_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17759__A _17759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22563_ _22146_/A _22558_/X _21826_/X _22562_/Y VGND VGND VPWR VPWR _22564_/A sky130_fd_sc_hd__a211o_4
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24302_ _25526_/CLK _17617_/X HRESETn VGND VGND VPWR VPWR _24302_/Q sky130_fd_sc_hd__dfrtp_4
X_21514_ _21284_/A VGND VGND VPWR VPWR _21514_/X sky130_fd_sc_hd__buf_2
X_25282_ _24252_/CLK _13701_/Y HRESETn VGND VGND VPWR VPWR _13693_/D sky130_fd_sc_hd__dfrtp_4
X_22494_ _14934_/Y _22442_/X _21573_/X _22493_/X VGND VGND VPWR VPWR _22494_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15724__A3 _15723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24233_ _23826_/CLK _18099_/X HRESETn VGND VGND VPWR VPWR _24233_/Q sky130_fd_sc_hd__dfrtp_4
X_21445_ _21196_/A VGND VGND VPWR VPWR _21469_/A sky130_fd_sc_hd__buf_2
XFILLER_119_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19974__A _19991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21376_ _21393_/A _20205_/Y VGND VGND VPWR VPWR _21376_/X sky130_fd_sc_hd__or2_4
XFILLER_134_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16134__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24164_ _24545_/CLK _18535_/X HRESETn VGND VGND VPWR VPWR _24164_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20327_ _20326_/Y VGND VGND VPWR VPWR _20327_/X sky130_fd_sc_hd__buf_2
X_23115_ _12277_/A _22980_/X _17742_/A _22906_/X VGND VGND VPWR VPWR _23115_/X sky130_fd_sc_hd__a2bb2o_4
X_24095_ _24097_/CLK _24095_/D HRESETn VGND VGND VPWR VPWR _12125_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_6_15_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20258_ _23434_/Q VGND VGND VPWR VPWR _20258_/Y sky130_fd_sc_hd__inv_2
X_23046_ _22769_/X _23042_/Y _22863_/X _23045_/X VGND VGND VPWR VPWR _23046_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20189_ _13748_/C _13752_/X _13735_/X _13762_/A VGND VGND VPWR VPWR _20189_/X sky130_fd_sc_hd__or4_4
XFILLER_62_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12431__A _12249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14999__B2 _16785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24997_ _24995_/CLK _24997_/D HRESETn VGND VGND VPWR VPWR _24997_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19387__B1 _19364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15660__A2 _15655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14750_ _14750_/A _14744_/X VGND VGND VPWR VPWR _14750_/X sky130_fd_sc_hd__and2_4
XFILLER_40_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11962_ _11650_/A _11959_/X _11702_/C _11961_/X VGND VGND VPWR VPWR _25489_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_1_1_1_HCLK clkbuf_1_1_0_HCLK/X VGND VGND VPWR VPWR clkbuf_2_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_23948_ _25199_/CLK _23948_/D HRESETn VGND VGND VPWR VPWR _23948_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21733__A2 _15708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13701_ _13701_/A VGND VGND VPWR VPWR _13701_/Y sky130_fd_sc_hd__inv_2
X_14681_ _14680_/X VGND VGND VPWR VPWR _14682_/B sky130_fd_sc_hd__buf_2
X_11893_ _11893_/A VGND VGND VPWR VPWR _11893_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23879_ _23869_/CLK _23879_/D VGND VGND VPWR VPWR _23879_/Q sky130_fd_sc_hd__dfxtp_4
X_16420_ _16418_/Y _16414_/X _16231_/X _16419_/X VGND VGND VPWR VPWR _16420_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24545__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13632_ _19014_/A _13631_/X _19014_/A _13631_/X VGND VGND VPWR VPWR _13633_/D sky130_fd_sc_hd__a2bb2o_4
X_16351_ _16349_/Y _16350_/X _16061_/X _16350_/X VGND VGND VPWR VPWR _24605_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21497__A1 _20333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13563_ _13562_/Y _25084_/Q _13562_/Y _25084_/Q VGND VGND VPWR VPWR _13564_/D sky130_fd_sc_hd__a2bb2o_4
X_15302_ _15422_/A VGND VGND VPWR VPWR _15388_/C sky130_fd_sc_hd__inv_2
XANTENNA__22294__B _22927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12514_ _12514_/A VGND VGND VPWR VPWR _12514_/Y sky130_fd_sc_hd__inv_2
X_19070_ _23857_/Q VGND VGND VPWR VPWR _19070_/Y sky130_fd_sc_hd__inv_2
X_16282_ _16282_/A VGND VGND VPWR VPWR _16282_/X sky130_fd_sc_hd__buf_2
X_13494_ _13493_/Y _13489_/X _13472_/X _13476_/Y VGND VGND VPWR VPWR _25304_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23238__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20095__A _20095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15715__A3 _15714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18021_ _18021_/A VGND VGND VPWR VPWR _18021_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15233_ _15233_/A _15233_/B VGND VGND VPWR VPWR _15235_/B sky130_fd_sc_hd__or2_4
X_12445_ _12199_/Y _12445_/B VGND VGND VPWR VPWR _12446_/C sky130_fd_sc_hd__nand2_4
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15164_ _15171_/B VGND VGND VPWR VPWR _15165_/B sky130_fd_sc_hd__buf_2
XANTENNA__21919__A _21944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12376_ _25350_/Q _12364_/Y _12363_/Y _24811_/Q VGND VGND VPWR VPWR _12380_/C sky130_fd_sc_hd__a2bb2o_4
X_14115_ _14115_/A _14115_/B _25205_/Q VGND VGND VPWR VPWR _14116_/B sky130_fd_sc_hd__or3_4
XFILLER_5_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15095_ _24982_/Q VGND VGND VPWR VPWR _15296_/A sky130_fd_sc_hd__inv_2
X_19972_ _17708_/A _18287_/A _18275_/A _19971_/X VGND VGND VPWR VPWR _19973_/A sky130_fd_sc_hd__or4_4
XFILLER_84_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25333__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14046_ _14045_/X VGND VGND VPWR VPWR _14046_/Y sky130_fd_sc_hd__inv_2
X_18923_ _19105_/A _17472_/A _18922_/X VGND VGND VPWR VPWR _18923_/X sky130_fd_sc_hd__or3_4
XFILLER_80_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18854_ _18854_/A _18854_/B _18852_/X _18853_/X VGND VGND VPWR VPWR _18865_/B sky130_fd_sc_hd__or4_4
XFILLER_95_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17805_ _17805_/A _17805_/B _17804_/X VGND VGND VPWR VPWR _17806_/A sky130_fd_sc_hd__or3_4
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17851__B _17846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15997_ _15996_/X VGND VGND VPWR VPWR _15997_/X sky130_fd_sc_hd__buf_2
X_18785_ _18678_/Y _18784_/X VGND VGND VPWR VPWR _18786_/D sky130_fd_sc_hd__or2_4
XANTENNA__22469__B _22468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14948_ _14947_/Y _24413_/Q _14947_/Y _24413_/Q VGND VGND VPWR VPWR _14951_/C sky130_fd_sc_hd__a2bb2o_4
X_17736_ _17700_/X _18319_/B _17734_/Y _21686_/A _17899_/A VGND VGND VPWR VPWR _24277_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21373__B _21373_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_35_0_HCLK clkbuf_8_34_0_HCLK/A VGND VGND VPWR VPWR _23818_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_63_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14879_ _14879_/A VGND VGND VPWR VPWR _14879_/Y sky130_fd_sc_hd__inv_2
X_17667_ _17676_/A _17676_/B VGND VGND VPWR VPWR _17674_/B sky130_fd_sc_hd__or2_4
Xclkbuf_8_98_0_HCLK clkbuf_8_99_0_HCLK/A VGND VGND VPWR VPWR _24356_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24286__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19406_ _18033_/B VGND VGND VPWR VPWR _19406_/Y sky130_fd_sc_hd__inv_2
X_16618_ _16618_/A VGND VGND VPWR VPWR _16618_/Y sky130_fd_sc_hd__inv_2
X_17598_ _17617_/A _17596_/X _17598_/C VGND VGND VPWR VPWR _24307_/D sky130_fd_sc_hd__and3_4
XANTENNA__18682__B _18682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16549_ _24531_/Q VGND VGND VPWR VPWR _16549_/Y sky130_fd_sc_hd__inv_2
X_19337_ _19336_/Y _19334_/X _19291_/X _19334_/X VGND VGND VPWR VPWR _19337_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22685__B1 _17755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19550__B1 _19389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19268_ _19268_/A VGND VGND VPWR VPWR _22205_/B sky130_fd_sc_hd__inv_2
XFILLER_31_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16364__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18219_ _17999_/A _18219_/B VGND VGND VPWR VPWR _18220_/C sky130_fd_sc_hd__or2_4
X_19199_ _19195_/Y _19198_/X _19155_/X _19198_/X VGND VGND VPWR VPWR _19199_/X sky130_fd_sc_hd__a2bb2o_4
X_21230_ _21372_/A VGND VGND VPWR VPWR _21253_/A sky130_fd_sc_hd__buf_2
XANTENNA__16116__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21161_ _17700_/C VGND VGND VPWR VPWR _21162_/A sky130_fd_sc_hd__inv_2
XFILLER_102_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17864__B1 _17790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21548__B _21548_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18203__A _18024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25074__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20112_ _20110_/Y _20106_/X _20085_/X _20111_/X VGND VGND VPWR VPWR _20112_/X sky130_fd_sc_hd__a2bb2o_4
X_21092_ _21029_/X _21090_/X _22664_/B _21091_/X VGND VGND VPWR VPWR _21093_/C sky130_fd_sc_hd__a211o_4
XANTENNA__25003__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20043_ _20043_/A _14697_/A _20043_/C _20043_/D VGND VGND VPWR VPWR _20044_/A sky130_fd_sc_hd__or4_4
XFILLER_86_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13347__A _13310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24920_ _25433_/CLK _24920_/D HRESETn VGND VGND VPWR VPWR _24920_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24851_ _25397_/CLK _15757_/X HRESETn VGND VGND VPWR VPWR _24851_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15562__A _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23802_ _23798_/CLK _23802_/D VGND VGND VPWR VPWR _13265_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_45_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24782_ _24800_/CLK _24782_/D HRESETn VGND VGND VPWR VPWR _22546_/A sky130_fd_sc_hd__dfrtp_4
X_21994_ _21994_/A VGND VGND VPWR VPWR _22727_/B sky130_fd_sc_hd__buf_2
XFILLER_96_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23733_ _23722_/CLK _19421_/X VGND VGND VPWR VPWR _19419_/A sky130_fd_sc_hd__dfxtp_4
X_20945_ _20818_/X _20944_/X _16648_/A _20864_/X VGND VGND VPWR VPWR _20945_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_6_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23664_ _23711_/CLK _19626_/X VGND VGND VPWR VPWR _19624_/A sky130_fd_sc_hd__dfxtp_4
X_20876_ _20860_/X _20875_/X _24479_/Q _20865_/X VGND VGND VPWR VPWR _20876_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25403_ _25400_/CLK _12689_/X HRESETn VGND VGND VPWR VPWR _25403_/Q sky130_fd_sc_hd__dfrtp_4
X_22615_ _24041_/Q _21302_/A _13132_/A _21304_/X VGND VGND VPWR VPWR _22615_/Y sky130_fd_sc_hd__a22oi_4
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16393__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23595_ _23434_/CLK _23595_/D VGND VGND VPWR VPWR _23595_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22140__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25334_ _25351_/CLK _25334_/D HRESETn VGND VGND VPWR VPWR _25334_/Q sky130_fd_sc_hd__dfrtp_4
X_22546_ _22546_/A _22587_/B VGND VGND VPWR VPWR _22546_/X sky130_fd_sc_hd__or2_4
XANTENNA__23938__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25265_ _25055_/CLK _13767_/X HRESETn VGND VGND VPWR VPWR _13757_/A sky130_fd_sc_hd__dfrtp_4
X_22477_ _21293_/A VGND VGND VPWR VPWR _22626_/B sky130_fd_sc_hd__buf_2
X_12230_ _25437_/Q _12228_/Y _12278_/B _22141_/A VGND VGND VPWR VPWR _12230_/X sky130_fd_sc_hd__a2bb2o_4
X_24216_ _24219_/CLK _18255_/X HRESETn VGND VGND VPWR VPWR _24216_/Q sky130_fd_sc_hd__dfrtp_4
X_21428_ _21323_/A VGND VGND VPWR VPWR _21428_/X sky130_fd_sc_hd__buf_2
XANTENNA__16107__B1 _15949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17718__A2_N _21465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25196_ _24942_/CLK _25196_/D HRESETn VGND VGND VPWR VPWR _20493_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22443__A3 _16728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12161_ _25153_/Q _12160_/X VGND VGND VPWR VPWR _12163_/A sky130_fd_sc_hd__or2_4
XANTENNA__16344__A2_N _16337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24147_ _24151_/CLK _18591_/X HRESETn VGND VGND VPWR VPWR _24147_/Q sky130_fd_sc_hd__dfrtp_4
X_21359_ _21351_/Y _21359_/B _21359_/C _21359_/D VGND VGND VPWR VPWR _21360_/B sky130_fd_sc_hd__and4_4
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18113__A _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12092_ _12092_/A VGND VGND VPWR VPWR _12092_/Y sky130_fd_sc_hd__inv_2
X_24078_ _24077_/CLK _24078_/D HRESETn VGND VGND VPWR VPWR _20428_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15920_ _15920_/A VGND VGND VPWR VPWR _15920_/Y sky130_fd_sc_hd__inv_2
X_23029_ _23024_/Y _23028_/Y _22850_/X VGND VGND VPWR VPWR _23030_/D sky130_fd_sc_hd__o21a_4
XFILLER_104_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21537__A1_N _17199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15851_ _21027_/A _15851_/B VGND VGND VPWR VPWR _15852_/A sky130_fd_sc_hd__or2_4
XANTENNA__24797__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14802_ _14802_/A _14802_/B _25039_/Q VGND VGND VPWR VPWR _14803_/B sky130_fd_sc_hd__or3_4
XANTENNA__24726__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15782_ _12050_/A _15782_/B _11716_/A _15991_/D VGND VGND VPWR VPWR _15782_/X sky130_fd_sc_hd__or4_4
X_18570_ _18555_/A _18566_/X _18570_/C VGND VGND VPWR VPWR _18570_/X sky130_fd_sc_hd__and3_4
XFILLER_40_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_251_0_HCLK clkbuf_7_125_0_HCLK/X VGND VGND VPWR VPWR _25397_/CLK sky130_fd_sc_hd__clkbuf_1
X_12994_ _25323_/Q VGND VGND VPWR VPWR _13106_/A sky130_fd_sc_hd__inv_2
X_14733_ _14732_/X VGND VGND VPWR VPWR _14733_/Y sky130_fd_sc_hd__inv_2
X_17521_ _24296_/Q VGND VGND VPWR VPWR _17521_/Y sky130_fd_sc_hd__inv_2
X_11945_ _19992_/A VGND VGND VPWR VPWR _19629_/A sky130_fd_sc_hd__buf_2
X_17452_ _24191_/Q _17452_/B VGND VGND VPWR VPWR _17453_/B sky130_fd_sc_hd__and2_4
XFILLER_32_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14664_ _14663_/X VGND VGND VPWR VPWR _18972_/A sky130_fd_sc_hd__buf_2
XANTENNA__15397__A1 _15073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11876_ _25499_/Q _11916_/A VGND VGND VPWR VPWR _11876_/X sky130_fd_sc_hd__and2_4
X_16403_ HWDATA[20] VGND VGND VPWR VPWR _16403_/X sky130_fd_sc_hd__buf_2
XANTENNA__15936__A3 HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13615_ _14645_/A VGND VGND VPWR VPWR _17995_/A sky130_fd_sc_hd__buf_2
X_17383_ _17344_/A _17377_/B _17383_/C VGND VGND VPWR VPWR _17383_/X sky130_fd_sc_hd__and3_4
XFILLER_38_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22667__B1 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14595_ _14592_/B _14586_/X _14594_/Y _14590_/X _13576_/A VGND VGND VPWR VPWR _14595_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22131__A2 _22122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16334_ _24611_/Q VGND VGND VPWR VPWR _16334_/Y sky130_fd_sc_hd__inv_2
X_19122_ _13402_/B VGND VGND VPWR VPWR _19122_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13546_ _25254_/Q VGND VGND VPWR VPWR _22612_/A sky130_fd_sc_hd__inv_2
XFILLER_41_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12080__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16346__B1 _16147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19053_ _19051_/Y _19052_/X _18961_/X _19052_/X VGND VGND VPWR VPWR _23863_/D sky130_fd_sc_hd__a2bb2o_4
X_16265_ _21322_/A VGND VGND VPWR VPWR _16265_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16453__D _11732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13477_ _13476_/Y VGND VGND VPWR VPWR _13477_/X sky130_fd_sc_hd__buf_2
XANTENNA__25514__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15216_ _15216_/A _15216_/B _15216_/C VGND VGND VPWR VPWR _15216_/X sky130_fd_sc_hd__and3_4
X_18004_ _18046_/A _18991_/A VGND VGND VPWR VPWR _18005_/C sky130_fd_sc_hd__or2_4
X_12428_ _12427_/X VGND VGND VPWR VPWR _25442_/D sky130_fd_sc_hd__inv_2
X_16196_ _16195_/Y _16193_/X _15942_/X _16193_/X VGND VGND VPWR VPWR _24662_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15147_ _15147_/A VGND VGND VPWR VPWR _15147_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15647__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12359_ _12358_/Y _24822_/Q _12358_/Y _24822_/Q VGND VGND VPWR VPWR _12359_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18023__A _14645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14551__A HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12183__A1_N _25426_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15078_ _24990_/Q VGND VGND VPWR VPWR _15331_/A sky130_fd_sc_hd__inv_2
X_19955_ _22245_/B _19952_/X _19615_/X _19952_/X VGND VGND VPWR VPWR _19955_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16484__A1_N _16483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14029_ _13997_/X _13998_/X _13990_/C _25221_/Q VGND VGND VPWR VPWR _14030_/B sky130_fd_sc_hd__a211o_4
X_18906_ _18906_/A VGND VGND VPWR VPWR _22062_/B sky130_fd_sc_hd__inv_2
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19886_ _21184_/B _19880_/X _19885_/X _19880_/A VGND VGND VPWR VPWR _19886_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13883__A1 _23989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_61_0_HCLK clkbuf_6_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18837_ _16535_/A _18633_/A _16535_/Y _18682_/B VGND VGND VPWR VPWR _18837_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16478__A _24558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24467__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18768_ _18768_/A _18765_/X VGND VGND VPWR VPWR _18768_/X sky130_fd_sc_hd__or2_4
XFILLER_97_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21158__B1 _16722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17719_ _24201_/Q VGND VGND VPWR VPWR _17719_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18699_ _18698_/X VGND VGND VPWR VPWR _18701_/B sky130_fd_sc_hd__inv_2
X_20730_ _20721_/X _20729_/X _24891_/Q _20726_/X VGND VGND VPWR VPWR _24008_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20661_ _14218_/Y _17404_/A _17387_/A _17401_/A VGND VGND VPWR VPWR _20662_/B sky130_fd_sc_hd__o22a_4
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22400_ _22400_/A _22266_/X VGND VGND VPWR VPWR _22400_/X sky130_fd_sc_hd__or2_4
XANTENNA__18433__A2_N _24168_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20592_ _20592_/A _20443_/B VGND VGND VPWR VPWR _20592_/Y sky130_fd_sc_hd__nand2_4
X_23380_ _24219_/CLK _20393_/X VGND VGND VPWR VPWR _21200_/A sky130_fd_sc_hd__dfxtp_4
X_22331_ _22327_/X _22330_/X _17722_/A VGND VGND VPWR VPWR _22331_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__25255__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25050_ _23494_/CLK _25050_/D HRESETn VGND VGND VPWR VPWR _14676_/A sky130_fd_sc_hd__dfrtp_4
X_22262_ _21270_/X _22224_/X _21950_/X _22261_/X VGND VGND VPWR VPWR _22263_/A sky130_fd_sc_hd__o22a_4
XANTENNA__18629__A2 _24142_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17756__B _17755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24001_ _24885_/CLK _20697_/Y HRESETn VGND VGND VPWR VPWR _13126_/A sky130_fd_sc_hd__dfrtp_4
X_21213_ _21069_/A VGND VGND VPWR VPWR _21859_/B sky130_fd_sc_hd__buf_2
XANTENNA__15557__A _16640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22193_ _21385_/A VGND VGND VPWR VPWR _22193_/X sky130_fd_sc_hd__buf_2
XFILLER_132_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21144_ _14214_/Y _14192_/A _21142_/Y _21143_/X VGND VGND VPWR VPWR _21144_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17772__A _16916_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21075_ _12983_/A _15654_/A _21031_/X _21074_/X VGND VGND VPWR VPWR _21075_/X sky130_fd_sc_hd__a211o_4
XFILLER_115_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20026_ _20026_/A VGND VGND VPWR VPWR _22253_/B sky130_fd_sc_hd__inv_2
XANTENNA__24890__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24903_ _24018_/CLK _15582_/X HRESETn VGND VGND VPWR VPWR _15579_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_74_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15292__A _15336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24834_ _24836_/CLK _24834_/D HRESETn VGND VGND VPWR VPWR _24834_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24137__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24765_ _24830_/CLK _15936_/X HRESETn VGND VGND VPWR VPWR _24765_/Q sky130_fd_sc_hd__dfrtp_4
X_21977_ _18359_/Y _21977_/B VGND VGND VPWR VPWR _21977_/X sky130_fd_sc_hd__and2_4
XFILLER_82_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19762__B1 _19715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11730_ _11730_/A _11730_/B _11730_/C _11730_/D VGND VGND VPWR VPWR _11731_/D sky130_fd_sc_hd__or4_4
XPHY_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23716_ _23683_/CLK _23716_/D VGND VGND VPWR VPWR _19466_/A sky130_fd_sc_hd__dfxtp_4
X_20928_ _20909_/X _20927_/X _24491_/Q _20913_/X VGND VGND VPWR VPWR _20928_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16576__B1 _16405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_81_0_HCLK clkbuf_8_81_0_HCLK/A VGND VGND VPWR VPWR _23964_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24696_ _24699_/CLK _16097_/X HRESETn VGND VGND VPWR VPWR _23219_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11661_ _24219_/Q VGND VGND VPWR VPWR _11661_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15016__A1_N _25022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23647_ _24288_/CLK _23647_/D VGND VGND VPWR VPWR _23647_/Q sky130_fd_sc_hd__dfxtp_4
X_20859_ _20858_/X VGND VGND VPWR VPWR _20859_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _13198_/X _13399_/X _25315_/Q _13258_/X VGND VGND VPWR VPWR _25315_/D sky130_fd_sc_hd__o22a_4
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14380_ _13976_/X _14380_/B VGND VGND VPWR VPWR _14380_/X sky130_fd_sc_hd__or2_4
XANTENNA__16328__B1 _16228_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12062__B1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20124__B2 _20105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23578_ _23545_/CLK _23578_/D VGND VGND VPWR VPWR _23578_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22853__A _22853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ _13428_/A _13329_/X _13330_/X VGND VGND VPWR VPWR _13331_/X sky130_fd_sc_hd__and3_4
XFILLER_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25317_ _25316_/CLK _25317_/D HRESETn VGND VGND VPWR VPWR _25317_/Q sky130_fd_sc_hd__dfrtp_4
X_22529_ _14900_/A _22523_/X _22524_/X _22528_/X VGND VGND VPWR VPWR _22530_/C sky130_fd_sc_hd__a211o_4
Xclkbuf_2_1_0_HCLK clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16050_ _16049_/Y _16047_/X _15897_/X _16047_/X VGND VGND VPWR VPWR _24713_/D sky130_fd_sc_hd__a2bb2o_4
X_13262_ _13212_/A VGND VGND VPWR VPWR _13402_/A sky130_fd_sc_hd__buf_2
XFILLER_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21469__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23074__B1 _21050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25248_ _25290_/CLK _13838_/X HRESETn VGND VGND VPWR VPWR _13551_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22416__A3 _22412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15001_ _15070_/B _24455_/Q _15070_/B _24455_/Q VGND VGND VPWR VPWR _15002_/D sky130_fd_sc_hd__a2bb2o_4
X_12213_ _12213_/A VGND VGND VPWR VPWR _12286_/C sky130_fd_sc_hd__inv_2
X_13193_ _13366_/A _13185_/X _13192_/X _11958_/X _11970_/C VGND VGND VPWR VPWR _13193_/X
+ sky130_fd_sc_hd__o32a_4
X_25179_ _25178_/CLK _14260_/X HRESETn VGND VGND VPWR VPWR _14254_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_29_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12144_ _25462_/Q _12143_/Y _25462_/Q _12143_/Y VGND VGND VPWR VPWR _12145_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24978__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16500__B1 _16325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19740_ _18254_/A VGND VGND VPWR VPWR _19740_/X sky130_fd_sc_hd__buf_2
XANTENNA__24907__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12075_ _12063_/Y _12074_/X _11833_/X _12074_/X VGND VGND VPWR VPWR _25473_/D sky130_fd_sc_hd__a2bb2o_4
X_16952_ _16932_/X _16952_/B _16952_/C _16952_/D VGND VGND VPWR VPWR _16952_/X sky130_fd_sc_hd__or4_4
XFILLER_110_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15903_ _12746_/Y _15900_/X _15623_/X _15900_/X VGND VGND VPWR VPWR _15903_/X sky130_fd_sc_hd__a2bb2o_4
X_19671_ _19671_/A VGND VGND VPWR VPWR _19671_/Y sky130_fd_sc_hd__inv_2
X_16883_ _20099_/A VGND VGND VPWR VPWR _19797_/A sky130_fd_sc_hd__buf_2
XANTENNA__20060__B1 _19797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24560__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18622_ _24526_/Q _24137_/Q _16562_/Y _18675_/A VGND VGND VPWR VPWR _18625_/C sky130_fd_sc_hd__o22a_4
XFILLER_66_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15834_ _12345_/Y _15833_/X _15627_/X _15833_/X VGND VGND VPWR VPWR _24812_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18553_ _18467_/A _18552_/Y VGND VGND VPWR VPWR _18553_/X sky130_fd_sc_hd__or2_4
X_12977_ _12979_/A _12970_/X _12977_/C VGND VGND VPWR VPWR _12977_/X sky130_fd_sc_hd__and3_4
X_15765_ _15742_/A VGND VGND VPWR VPWR _15765_/X sky130_fd_sc_hd__buf_2
XFILLER_45_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17504_ _11864_/Y _17577_/A _11864_/Y _17577_/A VGND VGND VPWR VPWR _17504_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15930__A _15795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11928_ _11928_/A VGND VGND VPWR VPWR _19615_/A sky130_fd_sc_hd__buf_2
X_14716_ _14716_/A VGND VGND VPWR VPWR _21633_/A sky130_fd_sc_hd__buf_2
X_15696_ _15687_/A _15687_/B _15695_/X VGND VGND VPWR VPWR _15696_/X sky130_fd_sc_hd__o21a_4
X_18484_ _24176_/Q _18483_/B VGND VGND VPWR VPWR _18484_/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14647_ _14646_/X VGND VGND VPWR VPWR _18005_/A sky130_fd_sc_hd__buf_2
X_17435_ _17434_/Y _17432_/X _16717_/X _17432_/X VGND VGND VPWR VPWR _17435_/X sky130_fd_sc_hd__a2bb2o_4
X_11859_ _11855_/Y _11848_/X _11858_/X _11848_/X VGND VGND VPWR VPWR _11859_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_109_0_HCLK clkbuf_7_54_0_HCLK/X VGND VGND VPWR VPWR _24033_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__19505__B1 _11948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22104__A2 _21009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13450__A _13450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ _25084_/Q _14577_/X _14575_/Y VGND VGND VPWR VPWR _14578_/X sky130_fd_sc_hd__o21a_4
X_17366_ _17369_/A _17369_/B VGND VGND VPWR VPWR _17370_/B sky130_fd_sc_hd__or2_4
XANTENNA__16319__B1 _15962_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19105_ _19105_/A _18331_/X _19683_/C VGND VGND VPWR VPWR _19106_/A sky130_fd_sc_hd__or3_4
X_13529_ _13529_/A VGND VGND VPWR VPWR _13529_/Y sky130_fd_sc_hd__inv_2
X_16317_ _16315_/Y _16311_/X _15959_/X _16316_/X VGND VGND VPWR VPWR _24618_/D sky130_fd_sc_hd__a2bb2o_4
X_17297_ _17266_/A _17295_/X _17296_/X VGND VGND VPWR VPWR _24353_/D sky130_fd_sc_hd__and3_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16761__A _24448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16248_ _16246_/Y _16241_/X _16143_/X _16247_/X VGND VGND VPWR VPWR _16248_/X sky130_fd_sc_hd__a2bb2o_4
X_19036_ _23868_/Q VGND VGND VPWR VPWR _19036_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17819__B1 _16955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16179_ _23323_/A VGND VGND VPWR VPWR _16179_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24648__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19938_ _19938_/A VGND VGND VPWR VPWR _19938_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18244__B1 _11821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19869_ _22328_/B _19868_/X _19612_/X _19868_/X VGND VGND VPWR VPWR _19869_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20051__B1 _19783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21900_ _21904_/A _20177_/Y VGND VGND VPWR VPWR _21901_/C sky130_fd_sc_hd__or2_4
XFILLER_95_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12518__A2_N _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22880_ _24552_/Q _22879_/X _22798_/X VGND VGND VPWR VPWR _22880_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16001__A _24732_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24230__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21831_ _14231_/Y _14223_/A _15470_/Y _15462_/A VGND VGND VPWR VPWR _21833_/B sky130_fd_sc_hd__o22a_4
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15840__A _14470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19744__B1 _19721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24550_ _24465_/CLK _16500_/X HRESETn VGND VGND VPWR VPWR _24550_/Q sky130_fd_sc_hd__dfrtp_4
X_21762_ _21618_/A _19920_/Y VGND VGND VPWR VPWR _21762_/X sky130_fd_sc_hd__or2_4
XANTENNA__21551__B1 _14868_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_68_0_HCLK clkbuf_7_69_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_68_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23501_ _24208_/CLK _20075_/X VGND VGND VPWR VPWR _23501_/Q sky130_fd_sc_hd__dfxtp_4
X_20713_ _20713_/A _20708_/Y VGND VGND VPWR VPWR _20713_/X sky130_fd_sc_hd__and2_4
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24481_ _24496_/CLK _16684_/X HRESETn VGND VGND VPWR VPWR _16682_/A sky130_fd_sc_hd__dfrtp_4
X_21693_ _23314_/B _21692_/X VGND VGND VPWR VPWR _21693_/X sky130_fd_sc_hd__and2_4
XANTENNA__25436__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12044__B1 _25475_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23432_ _23453_/CLK _23432_/D VGND VGND VPWR VPWR _23432_/Q sky130_fd_sc_hd__dfxtp_4
X_20644_ _14235_/Y _20628_/X _20619_/A _20643_/X VGND VGND VPWR VPWR _20645_/A sky130_fd_sc_hd__a211o_4
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23968__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23363_ _21006_/X VGND VGND VPWR VPWR IRQ[9] sky130_fd_sc_hd__buf_2
X_20575_ _18878_/X _20575_/B _20571_/C VGND VGND VPWR VPWR _20575_/X sky130_fd_sc_hd__and3_4
XANTENNA__16671__A _16664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25102_ _25178_/CLK _25102_/D HRESETn VGND VGND VPWR VPWR _25102_/Q sky130_fd_sc_hd__dfrtp_4
X_22314_ _21559_/X _22312_/X _21565_/X _22313_/X VGND VGND VPWR VPWR _22314_/X sky130_fd_sc_hd__o22a_4
X_23294_ _22701_/A _23291_/X _23294_/C VGND VGND VPWR VPWR _23299_/C sky130_fd_sc_hd__and3_4
X_25033_ _25029_/CLK _14860_/X HRESETn VGND VGND VPWR VPWR _14799_/C sky130_fd_sc_hd__dfrtp_4
X_22245_ _18293_/B _22245_/B VGND VGND VPWR VPWR _22247_/B sky130_fd_sc_hd__or2_4
XFILLER_117_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19982__A _19991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21082__A2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22176_ _22175_/X VGND VGND VPWR VPWR _22176_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24389__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21127_ _18894_/Y _21116_/Y _14377_/B _21126_/X VGND VGND VPWR VPWR _21127_/X sky130_fd_sc_hd__a211o_4
XFILLER_59_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24318__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21058_ _21029_/X _21056_/X _22664_/B _21057_/X VGND VGND VPWR VPWR _21059_/C sky130_fd_sc_hd__a211o_4
XFILLER_101_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15049__B1 _14888_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12900_ _12900_/A VGND VGND VPWR VPWR _12900_/Y sky130_fd_sc_hd__inv_2
X_20009_ _23529_/Q VGND VGND VPWR VPWR _21926_/B sky130_fd_sc_hd__inv_2
XFILLER_101_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13880_ _25232_/Q _13860_/X _21142_/A _13855_/X VGND VGND VPWR VPWR _13880_/X sky130_fd_sc_hd__o22a_4
XFILLER_98_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12831_ _12830_/Y _24802_/Q _12830_/Y _24802_/Q VGND VGND VPWR VPWR _12831_/X sky130_fd_sc_hd__a2bb2o_4
X_24817_ _24813_/CLK _24817_/D HRESETn VGND VGND VPWR VPWR _12305_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_41_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15550_ _15991_/A _15991_/B _15700_/C _15549_/X VGND VGND VPWR VPWR _15551_/B sky130_fd_sc_hd__or4_4
XANTENNA__19222__A _19221_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15750__A HWDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12762_ _12761_/Y _24772_/Q _12761_/Y _24772_/Q VGND VGND VPWR VPWR _12763_/D sky130_fd_sc_hd__a2bb2o_4
X_24748_ _24766_/CLK _15972_/X HRESETn VGND VGND VPWR VPWR _24748_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _20441_/A _20441_/B _14513_/A VGND VGND VPWR VPWR _14503_/B sky130_fd_sc_hd__or3_4
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _15640_/B VGND VGND VPWR VPWR _11719_/B sky130_fd_sc_hd__buf_2
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _14881_/Y _15476_/X _15480_/X _15476_/A VGND VGND VPWR VPWR _15481_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23953__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _12693_/B VGND VGND VPWR VPWR _12693_/X sky130_fd_sc_hd__or2_4
XFILLER_42_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24679_ _24334_/CLK _16139_/X HRESETn VGND VGND VPWR VPWR _22595_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _25124_/Q VGND VGND VPWR VPWR _22302_/A sky130_fd_sc_hd__inv_2
X_17220_ _22939_/A VGND VGND VPWR VPWR _17220_/Y sky130_fd_sc_hd__inv_2
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15772__A1 _15749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25106__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17151_ _17151_/A _17150_/X _17160_/C VGND VGND VPWR VPWR _24365_/D sky130_fd_sc_hd__and3_4
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ _14355_/X _14362_/X _25471_/Q _14360_/X VGND VGND VPWR VPWR _25146_/D sky130_fd_sc_hd__o22a_4
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16102_ _16100_/Y _16101_/X _11761_/X _16101_/X VGND VGND VPWR VPWR _16102_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13314_ _13314_/A _13309_/X _13313_/X VGND VGND VPWR VPWR _13315_/C sky130_fd_sc_hd__or3_4
X_17082_ _16976_/Y _17086_/B VGND VGND VPWR VPWR _17082_/Y sky130_fd_sc_hd__nand2_4
X_14294_ _14291_/C _14291_/D VGND VGND VPWR VPWR _14299_/A sky130_fd_sc_hd__or2_4
XANTENNA__16721__B1 _16720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16033_ _16033_/A VGND VGND VPWR VPWR _16033_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13535__B1 _13515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13245_ _13156_/X VGND VGND VPWR VPWR _13453_/A sky130_fd_sc_hd__buf_2
XFILLER_108_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13176_ _13143_/X _13163_/X _13175_/X VGND VGND VPWR VPWR _13176_/X sky130_fd_sc_hd__or3_4
XFILLER_83_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12127_ _12127_/A _12127_/B VGND VGND VPWR VPWR _12128_/B sky130_fd_sc_hd__and2_4
XANTENNA__24741__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17984_ _17975_/A VGND VGND VPWR VPWR _18168_/A sky130_fd_sc_hd__buf_2
XANTENNA__24059__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19723_ _23630_/Q VGND VGND VPWR VPWR _19723_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12058_ _19581_/B VGND VGND VPWR VPWR _15662_/B sky130_fd_sc_hd__buf_2
X_16935_ _16122_/Y _17826_/A _22976_/A _16900_/Y VGND VGND VPWR VPWR _16937_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11849__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24110__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19654_ _19652_/Y _19653_/X _19553_/X _19653_/X VGND VGND VPWR VPWR _19654_/X sky130_fd_sc_hd__a2bb2o_4
X_16866_ _16872_/A VGND VGND VPWR VPWR _16866_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16788__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18241__A3 _11812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22758__A _22725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18605_ _18598_/X _18600_/X _18602_/X _18605_/D VGND VGND VPWR VPWR _18605_/X sky130_fd_sc_hd__or4_4
X_15817_ _15817_/A VGND VGND VPWR VPWR _15817_/X sky130_fd_sc_hd__buf_2
X_19585_ _19585_/A VGND VGND VPWR VPWR _19586_/D sky130_fd_sc_hd__buf_2
XFILLER_18_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16797_ _16796_/X VGND VGND VPWR VPWR _16797_/X sky130_fd_sc_hd__buf_2
XFILLER_19_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18536_ _18461_/Y _18542_/B VGND VGND VPWR VPWR _18540_/B sky130_fd_sc_hd__or2_4
XFILLER_93_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15748_ _15728_/X _15742_/X _15747_/X _24855_/Q _15740_/X VGND VGND VPWR VPWR _24855_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_94_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18467_ _18467_/A VGND VGND VPWR VPWR _18467_/Y sky130_fd_sc_hd__inv_2
X_15679_ _24876_/Q VGND VGND VPWR VPWR _15682_/C sky130_fd_sc_hd__inv_2
XFILLER_34_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17418_ _16057_/A VGND VGND VPWR VPWR _17418_/X sky130_fd_sc_hd__buf_2
XFILLER_21_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18398_ _24155_/Q VGND VGND VPWR VPWR _18566_/A sky130_fd_sc_hd__inv_2
XANTENNA__12508__B _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12577__B2 _24857_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17349_ _17349_/A _17369_/A _17365_/A _17371_/A VGND VGND VPWR VPWR _17349_/X sky130_fd_sc_hd__or4_4
XANTENNA__21300__A3 _21296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20360_ _20360_/A VGND VGND VPWR VPWR _20360_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12329__B2 _12328_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19019_ _19012_/Y _19016_/X _19018_/X _19016_/X VGND VGND VPWR VPWR _19019_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24829__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20291_ _20289_/Y _20290_/X _19992_/X _20290_/X VGND VGND VPWR VPWR _20291_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22940__B _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22030_ _21664_/A _19894_/Y _21668_/A VGND VGND VPWR VPWR _22030_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22261__A1 _21260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21837__A _21837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15279__B1 _15174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24482__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24411__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23981_ _25219_/CLK _23981_/D HRESETn VGND VGND VPWR VPWR _17399_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_111_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12501__A1 _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_31_0_HCLK clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22932_ _23065_/A _22932_/B _22932_/C VGND VGND VPWR VPWR _22933_/D sky130_fd_sc_hd__and3_4
XFILLER_83_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16779__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22863_ _22186_/A VGND VGND VPWR VPWR _22863_/X sky130_fd_sc_hd__buf_2
XFILLER_71_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24602_ _24600_/CLK _24602_/D HRESETn VGND VGND VPWR VPWR _24602_/Q sky130_fd_sc_hd__dfrtp_4
X_21814_ _21681_/A _21806_/X _21814_/C VGND VGND VPWR VPWR _21814_/X sky130_fd_sc_hd__or3_4
XFILLER_58_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22794_ _22794_/A VGND VGND VPWR VPWR _22795_/A sky130_fd_sc_hd__inv_2
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24533_ _24561_/CLK _16546_/X HRESETn VGND VGND VPWR VPWR _16541_/A sky130_fd_sc_hd__dfrtp_4
X_21745_ _21596_/A _21745_/B VGND VGND VPWR VPWR _21747_/B sky130_fd_sc_hd__or2_4
XFILLER_12_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25270__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24473__CLK _24581_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24464_ _25001_/CLK _16731_/X HRESETn VGND VGND VPWR VPWR _24464_/Q sky130_fd_sc_hd__dfrtp_4
X_21676_ _21650_/A _19573_/Y VGND VGND VPWR VPWR _21676_/X sky130_fd_sc_hd__or2_4
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12568__B2 _24856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23415_ _23714_/CLK _20309_/X VGND VGND VPWR VPWR _20308_/A sky130_fd_sc_hd__dfxtp_4
X_20627_ _20627_/A VGND VGND VPWR VPWR _20627_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_155_0_HCLK clkbuf_7_77_0_HCLK/X VGND VGND VPWR VPWR _24285_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24395_ _23846_/CLK _16882_/X HRESETn VGND VGND VPWR VPWR _20096_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23346_ VGND VGND VPWR VPWR _23346_/HI IRQ[12] sky130_fd_sc_hd__conb_1
X_20558_ _18875_/B _20557_/Y _20558_/C VGND VGND VPWR VPWR _20558_/X sky130_fd_sc_hd__and3_4
XANTENNA__16703__B1 _16521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23277_ _23276_/X VGND VGND VPWR VPWR _23277_/Y sky130_fd_sc_hd__inv_2
X_20489_ _14205_/A _20487_/X _20481_/C _20488_/X VGND VGND VPWR VPWR _20489_/Y sky130_fd_sc_hd__a22oi_4
X_13030_ _13030_/A _13038_/B VGND VGND VPWR VPWR _13035_/B sky130_fd_sc_hd__or2_4
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25016_ _25016_/CLK _15216_/X HRESETn VGND VGND VPWR VPWR _15065_/A sky130_fd_sc_hd__dfrtp_4
X_22228_ _21668_/A _22226_/X _22227_/X VGND VGND VPWR VPWR _22228_/X sky130_fd_sc_hd__and3_4
XFILLER_121_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15745__A HWDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22159_ _14439_/Y _21352_/A _14456_/Y _21355_/A VGND VGND VPWR VPWR _22159_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14981_ _14975_/Y VGND VGND VPWR VPWR _14981_/X sky130_fd_sc_hd__buf_2
XFILLER_82_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20015__B1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14493__B2 _14481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16720_ _16720_/A VGND VGND VPWR VPWR _16720_/X sky130_fd_sc_hd__buf_2
X_13932_ _24961_/Q VGND VGND VPWR VPWR _13932_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13863_ _13850_/Y VGND VGND VPWR VPWR _13863_/X sky130_fd_sc_hd__buf_2
X_16651_ _16658_/A VGND VGND VPWR VPWR _16651_/X sky130_fd_sc_hd__buf_2
XANTENNA__25358__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12814_ _12927_/A _24787_/Q _12927_/A _24787_/Q VGND VGND VPWR VPWR _12814_/X sky130_fd_sc_hd__a2bb2o_4
X_15602_ _24894_/Q VGND VGND VPWR VPWR _15602_/Y sky130_fd_sc_hd__inv_2
X_19370_ _11856_/X VGND VGND VPWR VPWR _19370_/X sky130_fd_sc_hd__buf_2
X_13794_ _21498_/A VGND VGND VPWR VPWR _13795_/D sky130_fd_sc_hd__buf_2
X_16582_ _16550_/A VGND VGND VPWR VPWR _16583_/A sky130_fd_sc_hd__buf_2
XANTENNA__21515__B1 _25509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18321_ _24198_/Q _18320_/Y _17891_/Y VGND VGND VPWR VPWR _24198_/D sky130_fd_sc_hd__o21a_4
X_12745_ _12744_/Y _24803_/Q _12744_/Y _24803_/Q VGND VGND VPWR VPWR _12745_/X sky130_fd_sc_hd__a2bb2o_4
X_15533_ _15662_/A VGND VGND VPWR VPWR _15533_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14096__A scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_51_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15464_ _15461_/Y _15463_/X _14411_/X _15463_/X VGND VGND VPWR VPWR _24945_/D sky130_fd_sc_hd__a2bb2o_4
X_18252_ _18235_/X _18237_/X _15836_/X _21967_/A _18238_/X VGND VGND VPWR VPWR _24217_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_124_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12676_ _12681_/A _12683_/A _12679_/A _12689_/B VGND VGND VPWR VPWR _12682_/B sky130_fd_sc_hd__or4_4
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _14128_/Y _14409_/X _14414_/X _14409_/X VGND VGND VPWR VPWR _25131_/D sky130_fd_sc_hd__a2bb2o_4
X_17203_ _22815_/A VGND VGND VPWR VPWR _17203_/Y sky130_fd_sc_hd__inv_2
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21818__A1 _21636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15395_ _15301_/D _15398_/B VGND VGND VPWR VPWR _15399_/B sky130_fd_sc_hd__or2_4
X_18183_ _18215_/A _19007_/A VGND VGND VPWR VPWR _18184_/C sky130_fd_sc_hd__or2_4
XFILLER_50_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ _14337_/Y _14345_/X _14325_/X VGND VGND VPWR VPWR _14346_/Y sky130_fd_sc_hd__a21oi_4
X_17134_ _17038_/A _17134_/B VGND VGND VPWR VPWR _17135_/B sky130_fd_sc_hd__or2_4
XFILLER_11_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24993__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17498__B2 _24294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22491__B2 _22288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13508__B1 _11847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17065_ _17050_/A _17260_/A VGND VGND VPWR VPWR _17065_/X sky130_fd_sc_hd__and2_4
XANTENNA__24922__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14277_ _14249_/A VGND VGND VPWR VPWR _14278_/A sky130_fd_sc_hd__inv_2
XANTENNA__16170__A1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12344__A _24808_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16016_ _16014_/Y _16010_/X _15949_/X _16015_/X VGND VGND VPWR VPWR _24727_/D sky130_fd_sc_hd__a2bb2o_4
X_13228_ _13417_/A _23507_/Q VGND VGND VPWR VPWR _13229_/C sky130_fd_sc_hd__or2_4
XFILLER_124_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21657__A _21465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_14_0_HCLK_A clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13159_ _13180_/A _13159_/B VGND VGND VPWR VPWR _13159_/X sky130_fd_sc_hd__or2_4
XFILLER_135_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17967_ _18024_/A _17967_/B VGND VGND VPWR VPWR _17967_/X sky130_fd_sc_hd__or2_4
XFILLER_61_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19706_ _19705_/X VGND VGND VPWR VPWR _19706_/Y sky130_fd_sc_hd__inv_2
X_16918_ _16918_/A VGND VGND VPWR VPWR _16918_/Y sky130_fd_sc_hd__inv_2
X_17898_ _17897_/X VGND VGND VPWR VPWR _17898_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19637_ _18333_/X _18334_/X _19728_/A _19683_/B VGND VGND VPWR VPWR _19638_/A sky130_fd_sc_hd__or4_4
X_16849_ _16847_/Y _16844_/X _16782_/X _16848_/X VGND VGND VPWR VPWR _24405_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21823__C _21784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25099__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19568_ _22023_/B _19562_/X _11939_/X _19567_/X VGND VGND VPWR VPWR _23682_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25028__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18519_ _18821_/B _18519_/B _18518_/X VGND VGND VPWR VPWR _18520_/A sky130_fd_sc_hd__or3_4
X_19499_ _23706_/Q VGND VGND VPWR VPWR _22004_/B sky130_fd_sc_hd__inv_2
XANTENNA__25117__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21521__A3 _21514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21530_ _22464_/A VGND VGND VPWR VPWR _21530_/X sky130_fd_sc_hd__buf_2
XFILLER_90_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11744__A1_N _11706_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21461_ _21452_/X _21460_/X _17722_/X VGND VGND VPWR VPWR _21461_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_8_228_0_HCLK clkbuf_8_229_0_HCLK/A VGND VGND VPWR VPWR _24766_/CLK sky130_fd_sc_hd__clkbuf_1
X_23200_ _23200_/A _23057_/X VGND VGND VPWR VPWR _23203_/B sky130_fd_sc_hd__or2_4
X_20412_ _20399_/Y VGND VGND VPWR VPWR _20412_/X sky130_fd_sc_hd__buf_2
XFILLER_105_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24180_ _23933_/CLK _24180_/D HRESETn VGND VGND VPWR VPWR _18383_/A sky130_fd_sc_hd__dfrtp_4
X_21392_ _21371_/A _19861_/Y VGND VGND VPWR VPWR _21392_/X sky130_fd_sc_hd__or2_4
XANTENNA__24663__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23131_ _16476_/A _22879_/X _23130_/X VGND VGND VPWR VPWR _23131_/X sky130_fd_sc_hd__o21a_4
X_20343_ _20342_/Y _20340_/X _19615_/A _20340_/X VGND VGND VPWR VPWR _23402_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12254__A _25424_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23062_ _24590_/Q _23171_/B VGND VGND VPWR VPWR _23065_/B sky130_fd_sc_hd__or2_4
X_20274_ _23428_/Q _20273_/Y _23968_/D _20272_/X VGND VGND VPWR VPWR _20274_/X sky130_fd_sc_hd__o22a_4
X_22013_ _22016_/A _22013_/B VGND VGND VPWR VPWR _22015_/B sky130_fd_sc_hd__or2_4
XFILLER_102_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12701__B _12665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22537__A2 _22533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23964_ _23964_/CLK _23964_/D HRESETn VGND VGND VPWR VPWR _23964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22915_ _22915_/A VGND VGND VPWR VPWR _23052_/B sky130_fd_sc_hd__buf_2
XFILLER_56_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23895_ _23905_/CLK _23895_/D VGND VGND VPWR VPWR _18959_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__15424__B1 _15318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25451__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22846_ _22836_/B VGND VGND VPWR VPWR _22846_/X sky130_fd_sc_hd__buf_2
XANTENNA__12789__A1 _25357_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22777_ _22769_/X _22773_/Y _22483_/X _22776_/X VGND VGND VPWR VPWR _22777_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _12529_/Y _24842_/Q _12529_/Y _24842_/Q VGND VGND VPWR VPWR _12530_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_6_38_0_HCLK clkbuf_5_19_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_38_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24516_ _24517_/CLK _24516_/D HRESETn VGND VGND VPWR VPWR _16587_/A sky130_fd_sc_hd__dfrtp_4
X_21728_ _21547_/Y _21721_/X _21723_/X _21727_/Y VGND VGND VPWR VPWR _21744_/B sky130_fd_sc_hd__a211o_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25496_ _25497_/CLK _11931_/X HRESETn VGND VGND VPWR VPWR _11928_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12461_ _12461_/A VGND VGND VPWR VPWR _12461_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24447_ _24447_/CLK _24447_/D HRESETn VGND VGND VPWR VPWR _24447_/Q sky130_fd_sc_hd__dfrtp_4
X_21659_ _21467_/A _21659_/B _21659_/C VGND VGND VPWR VPWR _21659_/X sky130_fd_sc_hd__and3_4
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14200_ _14200_/A VGND VGND VPWR VPWR _14201_/A sky130_fd_sc_hd__buf_2
XANTENNA__17020__A _17260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15180_ _15180_/A _15180_/B VGND VGND VPWR VPWR _15181_/C sky130_fd_sc_hd__or2_4
X_12392_ _12385_/A _12385_/B _12391_/X VGND VGND VPWR VPWR _12392_/X sky130_fd_sc_hd__or3_4
XFILLER_137_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24378_ _24720_/CLK _24378_/D HRESETn VGND VGND VPWR VPWR _16987_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14131_ _14125_/X _14130_/X _14097_/A _14125_/X VGND VGND VPWR VPWR _25211_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_14_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23329_ _24432_/Q _22135_/X _22797_/X _23328_/X VGND VGND VPWR VPWR _23330_/C sky130_fd_sc_hd__a211o_4
XFILLER_125_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24333__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14062_ _13976_/X VGND VGND VPWR VPWR _20452_/B sky130_fd_sc_hd__inv_2
XANTENNA__18429__B1 _16237_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14163__B1 _25121_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13013_ _13013_/A VGND VGND VPWR VPWR _13013_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20236__B1 _19755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18870_ _20537_/A _20537_/B VGND VGND VPWR VPWR _20539_/A sky130_fd_sc_hd__or2_4
X_17821_ _17758_/D _17818_/D VGND VGND VPWR VPWR _17825_/A sky130_fd_sc_hd__or2_4
XANTENNA__22528__A2 _22525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25539__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17752_ _17752_/A VGND VGND VPWR VPWR _17759_/A sky130_fd_sc_hd__inv_2
X_14964_ _25017_/Q VGND VGND VPWR VPWR _15000_/A sky130_fd_sc_hd__inv_2
XANTENNA__21736__B1 _22444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16703_ _16702_/Y _16700_/X _16521_/X _16700_/X VGND VGND VPWR VPWR _24473_/D sky130_fd_sc_hd__a2bb2o_4
X_13915_ _13945_/A _13913_/Y _13893_/B _13914_/X VGND VGND VPWR VPWR _13916_/A sky130_fd_sc_hd__or4_4
XFILLER_48_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17504__A1_N _11864_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17683_ _17683_/A VGND VGND VPWR VPWR _17683_/Y sky130_fd_sc_hd__inv_2
X_14895_ _15197_/A _16809_/A _14893_/Y _16809_/A VGND VGND VPWR VPWR _14895_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19422_ _17953_/B VGND VGND VPWR VPWR _19422_/Y sky130_fd_sc_hd__inv_2
X_16634_ _16630_/Y _16634_/B VGND VGND VPWR VPWR _16634_/X sky130_fd_sc_hd__or2_4
XFILLER_74_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13846_ _13846_/A VGND VGND VPWR VPWR _21368_/A sky130_fd_sc_hd__inv_2
XFILLER_63_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19353_ _17945_/B VGND VGND VPWR VPWR _19353_/Y sky130_fd_sc_hd__inv_2
X_13777_ _13777_/A VGND VGND VPWR VPWR _14406_/A sky130_fd_sc_hd__buf_2
X_16565_ _24525_/Q VGND VGND VPWR VPWR _16565_/Y sky130_fd_sc_hd__inv_2
X_18304_ _18301_/X VGND VGND VPWR VPWR _18304_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22700__A2 _22406_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15516_ _15516_/A VGND VGND VPWR VPWR _15535_/A sky130_fd_sc_hd__buf_2
X_12728_ _12728_/A _12735_/A VGND VGND VPWR VPWR _12737_/A sky130_fd_sc_hd__or2_4
X_19284_ _13158_/B VGND VGND VPWR VPWR _19284_/Y sky130_fd_sc_hd__inv_2
X_16496_ _16495_/Y _16491_/X _16410_/X _16491_/X VGND VGND VPWR VPWR _16496_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18235_ _18235_/A VGND VGND VPWR VPWR _18235_/X sky130_fd_sc_hd__buf_2
X_12659_ _12659_/A _12659_/B VGND VGND VPWR VPWR _12660_/C sky130_fd_sc_hd__or2_4
X_15447_ _13889_/C _15437_/X _15446_/X _13920_/X _15444_/X VGND VGND VPWR VPWR _15447_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18166_ _18023_/X _18164_/X _18165_/X VGND VGND VPWR VPWR _18166_/X sky130_fd_sc_hd__and3_4
X_15378_ _15285_/X VGND VGND VPWR VPWR _15384_/A sky130_fd_sc_hd__buf_2
XANTENNA__22771__A _24615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17117_ _17116_/X VGND VGND VPWR VPWR _17117_/Y sky130_fd_sc_hd__inv_2
X_14329_ _14329_/A _24094_/Q VGND VGND VPWR VPWR _14330_/A sky130_fd_sc_hd__or2_4
X_18097_ _18097_/A _18097_/B _18096_/X VGND VGND VPWR VPWR _18097_/X sky130_fd_sc_hd__and3_4
XFILLER_128_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24074__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_58_0_HCLK clkbuf_8_59_0_HCLK/A VGND VGND VPWR VPWR _24219_/CLK sky130_fd_sc_hd__clkbuf_1
X_17048_ _17048_/A _17048_/B _17029_/X _17048_/D VGND VGND VPWR VPWR _17066_/B sky130_fd_sc_hd__or4_4
XANTENNA__20227__B1 _18267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24003__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20778__B2 _20774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18999_ _18995_/Y _18989_/X _18997_/X _18998_/X VGND VGND VPWR VPWR _23882_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23177__C1 _23176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23107__A _24624_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20961_ _12134_/A _12159_/X VGND VGND VPWR VPWR _20961_/X sky130_fd_sc_hd__and2_4
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22700_ _16587_/A _22406_/B _21556_/X _22699_/X VGND VGND VPWR VPWR _22701_/C sky130_fd_sc_hd__a211o_4
XANTENNA__13633__A _13634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23680_ _24930_/CLK _23680_/D VGND VGND VPWR VPWR _23680_/Q sky130_fd_sc_hd__dfxtp_4
X_20892_ _24046_/Q VGND VGND VPWR VPWR _20892_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21272__D _21272_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22631_ _22631_/A _23035_/A VGND VGND VPWR VPWR _22631_/X sky130_fd_sc_hd__or2_4
XFILLER_41_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22152__B1 _22997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25350_ _25351_/CLK _25350_/D HRESETn VGND VGND VPWR VPWR _25350_/Q sky130_fd_sc_hd__dfrtp_4
X_22562_ _21580_/A _22562_/B VGND VGND VPWR VPWR _22562_/Y sky130_fd_sc_hd__nor2_4
XFILLER_70_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24301_ _25436_/CLK _17620_/X HRESETn VGND VGND VPWR VPWR _24301_/Q sky130_fd_sc_hd__dfrtp_4
X_21513_ _21513_/A _22998_/A VGND VGND VPWR VPWR _21513_/X sky130_fd_sc_hd__or2_4
XFILLER_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24844__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25281_ _24252_/CLK _13704_/X HRESETn VGND VGND VPWR VPWR _13693_/C sky130_fd_sc_hd__dfrtp_4
X_22493_ _15013_/Y _22493_/B VGND VGND VPWR VPWR _22493_/X sky130_fd_sc_hd__and2_4
XFILLER_72_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24232_ _23826_/CLK _24232_/D HRESETn VGND VGND VPWR VPWR _24232_/Q sky130_fd_sc_hd__dfrtp_4
X_21444_ _21444_/A VGND VGND VPWR VPWR _21510_/C sky130_fd_sc_hd__inv_2
XFILLER_124_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24163_ _24545_/CLK _18539_/X HRESETn VGND VGND VPWR VPWR _18420_/A sky130_fd_sc_hd__dfrtp_4
X_21375_ _21371_/A _21375_/B VGND VGND VPWR VPWR _21377_/B sky130_fd_sc_hd__or2_4
XFILLER_134_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23114_ _23114_/A _23114_/B _23104_/X _23113_/X VGND VGND VPWR VPWR _23114_/X sky130_fd_sc_hd__or4_4
X_20326_ _20326_/A VGND VGND VPWR VPWR _20326_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21297__A _21314_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24094_ _24102_/CLK _14331_/Y HRESETn VGND VGND VPWR VPWR _24094_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20218__B1 _19758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15893__B1 _22623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23045_ _22975_/X _23043_/X _23044_/X _25530_/Q _22775_/X VGND VGND VPWR VPWR _23045_/X
+ sky130_fd_sc_hd__a32o_4
X_20257_ _22189_/B _20254_/X _19780_/A _20254_/X VGND VGND VPWR VPWR _20257_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20769__B2 _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18831__B1 _16533_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20188_ _23460_/Q VGND VGND VPWR VPWR _22357_/B sky130_fd_sc_hd__inv_2
XFILLER_89_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12431__B _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24996_ _24995_/CLK _24996_/D HRESETn VGND VGND VPWR VPWR _14990_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11961_ _11961_/A _11967_/D _11647_/X _11967_/B VGND VGND VPWR VPWR _11961_/X sky130_fd_sc_hd__and4_4
XANTENNA__15660__A3 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23947_ _25098_/CLK sda_i_S4 HRESETn VGND VGND VPWR VPWR _23948_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13700_ _11673_/Y _13695_/X _13699_/X _13695_/B VGND VGND VPWR VPWR _13701_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22930__A2 _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14680_ _21371_/A VGND VGND VPWR VPWR _14680_/X sky130_fd_sc_hd__buf_2
X_11892_ _11892_/A _11887_/X VGND VGND VPWR VPWR _11893_/A sky130_fd_sc_hd__or2_4
X_23878_ _23869_/CLK _23878_/D VGND VGND VPWR VPWR _19007_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16070__B1 _15474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13631_ _18079_/A _13605_/X _17928_/A _13606_/Y VGND VGND VPWR VPWR _13631_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22829_ _23126_/A _22825_/X _22826_/X _22828_/X VGND VGND VPWR VPWR _22830_/A sky130_fd_sc_hd__o22a_4
XFILLER_71_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13562_ _25256_/Q VGND VGND VPWR VPWR _13562_/Y sky130_fd_sc_hd__inv_2
X_16350_ _16324_/A VGND VGND VPWR VPWR _16350_/X sky130_fd_sc_hd__buf_2
XFILLER_125_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12513_ _12512_/Y _24873_/Q _12512_/Y _24873_/Q VGND VGND VPWR VPWR _12513_/X sky130_fd_sc_hd__a2bb2o_4
X_15301_ _15159_/X _15388_/B _15073_/Y _15301_/D VGND VGND VPWR VPWR _15301_/X sky130_fd_sc_hd__or4_4
X_16281_ _16280_/X VGND VGND VPWR VPWR _16282_/A sky130_fd_sc_hd__buf_2
XANTENNA__24585__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13493_ _25304_/Q VGND VGND VPWR VPWR _13493_/Y sky130_fd_sc_hd__inv_2
X_25479_ _25284_/CLK _25479_/D HRESETn VGND VGND VPWR VPWR _12036_/A sky130_fd_sc_hd__dfrtp_4
X_18020_ _15695_/X _17994_/X _18018_/X _24236_/Q _18019_/X VGND VGND VPWR VPWR _18020_/X
+ sky130_fd_sc_hd__o32a_4
X_12444_ _12286_/B _12447_/A VGND VGND VPWR VPWR _12445_/B sky130_fd_sc_hd__or2_4
X_15232_ _15232_/A VGND VGND VPWR VPWR _15233_/B sky130_fd_sc_hd__inv_2
XANTENNA__24514__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14923__A2 _14922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12395__C1 _12394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_211_0_HCLK clkbuf_8_211_0_HCLK/A VGND VGND VPWR VPWR _24407_/CLK sky130_fd_sc_hd__clkbuf_1
X_15163_ _15121_/X _15162_/X VGND VGND VPWR VPWR _15171_/B sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_3_0_0_HCLK_A clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12375_ _12374_/Y _24837_/Q _12374_/Y _24837_/Q VGND VGND VPWR VPWR _12380_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14114_ _14099_/C _14113_/X _14100_/A VGND VGND VPWR VPWR _14115_/B sky130_fd_sc_hd__or3_4
X_15094_ _15085_/X _15088_/X _15091_/X _15093_/X VGND VGND VPWR VPWR _15121_/B sky130_fd_sc_hd__or4_4
X_19971_ _24205_/Q VGND VGND VPWR VPWR _19971_/X sky130_fd_sc_hd__buf_2
XANTENNA__15884__B1 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14045_ _14045_/A _14045_/B _14025_/C _13992_/X VGND VGND VPWR VPWR _14045_/X sky130_fd_sc_hd__or4_4
X_18922_ _17466_/Y _19219_/C _17459_/X VGND VGND VPWR VPWR _18922_/X sky130_fd_sc_hd__or3_4
XFILLER_122_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18853_ _16508_/Y _18686_/A _16508_/Y _18686_/A VGND VGND VPWR VPWR _18853_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21935__A _21458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21705__A1_N _17244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25373__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17804_ _17792_/B _17771_/B _16943_/Y VGND VGND VPWR VPWR _17804_/X sky130_fd_sc_hd__o21a_4
XFILLER_79_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18784_ _18683_/D _18783_/X VGND VGND VPWR VPWR _18784_/X sky130_fd_sc_hd__or2_4
X_15996_ _15995_/X VGND VGND VPWR VPWR _15996_/X sky130_fd_sc_hd__buf_2
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17851__C _16898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12060__C _15652_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25302__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17735_ _17700_/X _17735_/B _24198_/Q VGND VGND VPWR VPWR _17899_/A sky130_fd_sc_hd__or3_4
XANTENNA__15651__A3 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14947_ _14947_/A VGND VGND VPWR VPWR _14947_/Y sky130_fd_sc_hd__inv_2
X_17666_ _17512_/Y _17665_/X VGND VGND VPWR VPWR _17676_/B sky130_fd_sc_hd__or2_4
X_14878_ _14876_/Y _14810_/X _14835_/X _14877_/Y VGND VGND VPWR VPWR _14879_/A sky130_fd_sc_hd__o22a_4
XFILLER_1_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22766__A _21418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19405_ _19403_/Y _19401_/X _19404_/X _19401_/X VGND VGND VPWR VPWR _19405_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16617_ _16616_/Y _16614_/X _16359_/X _16614_/X VGND VGND VPWR VPWR _16617_/X sky130_fd_sc_hd__a2bb2o_4
X_13829_ _13822_/A VGND VGND VPWR VPWR _13829_/X sky130_fd_sc_hd__buf_2
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17597_ _17597_/A _17597_/B VGND VGND VPWR VPWR _17598_/C sky130_fd_sc_hd__or2_4
XFILLER_16_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22134__B1 _22792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19336_ _18002_/B VGND VGND VPWR VPWR _19336_/Y sky130_fd_sc_hd__inv_2
X_16548_ _16547_/Y _16545_/X _16285_/X _16545_/X VGND VGND VPWR VPWR _16548_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22685__A1 _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_21_0_HCLK clkbuf_6_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_42_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19267_ _19262_/Y _19266_/X _16863_/X _19266_/X VGND VGND VPWR VPWR _19267_/X sky130_fd_sc_hd__a2bb2o_4
X_16479_ _16474_/A VGND VGND VPWR VPWR _16479_/X sky130_fd_sc_hd__buf_2
X_18218_ _18186_/A _23829_/Q VGND VGND VPWR VPWR _18218_/X sky130_fd_sc_hd__or2_4
XANTENNA__24255__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19198_ _19197_/X VGND VGND VPWR VPWR _19198_/X sky130_fd_sc_hd__buf_2
XFILLER_102_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18149_ _18000_/A _18149_/B _18149_/C VGND VGND VPWR VPWR _18153_/B sky130_fd_sc_hd__and3_4
XANTENNA__20999__A1 _23962_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21160_ _17447_/X VGND VGND VPWR VPWR _21160_/X sky130_fd_sc_hd__buf_2
XANTENNA__17864__A1 _17846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20111_ _20105_/X VGND VGND VPWR VPWR _20111_/X sky130_fd_sc_hd__buf_2
XANTENNA__20914__A1_N _20909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19066__B1 _18993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21091_ _21091_/A _21038_/B VGND VGND VPWR VPWR _21091_/X sky130_fd_sc_hd__and2_4
XFILLER_63_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20042_ _20042_/A VGND VGND VPWR VPWR _22368_/B sky130_fd_sc_hd__inv_2
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15890__A3 _11800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24850_ _25397_/CLK _15760_/X HRESETn VGND VGND VPWR VPWR _24850_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14992__A2_N _24434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25043__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23801_ _23798_/CLK _23801_/D VGND VGND VPWR VPWR _13303_/B sky130_fd_sc_hd__dfxtp_4
X_24781_ _24813_/CLK _15899_/X HRESETn VGND VGND VPWR VPWR _24781_/Q sky130_fd_sc_hd__dfrtp_4
X_21993_ _13784_/D _23340_/B VGND VGND VPWR VPWR _21993_/Y sky130_fd_sc_hd__nand2_4
X_23732_ _23722_/CLK _23732_/D VGND VGND VPWR VPWR _17953_/B sky130_fd_sc_hd__dfxtp_4
X_20944_ _20942_/Y _20939_/X _20943_/X VGND VGND VPWR VPWR _20944_/X sky130_fd_sc_hd__o21a_4
XFILLER_22_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_103_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_207_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ _23398_/CLK _19630_/X VGND VGND VPWR VPWR _19627_/A sky130_fd_sc_hd__dfxtp_4
X_20875_ _20873_/Y _20870_/Y _20879_/B VGND VGND VPWR VPWR _20875_/X sky130_fd_sc_hd__o21a_4
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22395__B _21026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25402_ _25400_/CLK _12691_/Y HRESETn VGND VGND VPWR VPWR _12567_/A sky130_fd_sc_hd__dfrtp_4
X_22614_ _22505_/X _22612_/X _21950_/X _22613_/Y VGND VGND VPWR VPWR _22614_/X sky130_fd_sc_hd__o22a_4
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23594_ _23562_/CLK _23594_/D VGND VGND VPWR VPWR _19828_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25333_ _25351_/CLK _13089_/X HRESETn VGND VGND VPWR VPWR _25333_/Q sky130_fd_sc_hd__dfrtp_4
X_22545_ _22544_/X VGND VGND VPWR VPWR _22545_/X sky130_fd_sc_hd__buf_2
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25264_ _25264_/CLK _25264_/D HRESETn VGND VGND VPWR VPWR _13757_/B sky130_fd_sc_hd__dfrtp_4
X_22476_ _21511_/X VGND VGND VPWR VPWR _22476_/X sky130_fd_sc_hd__buf_2
XFILLER_136_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16605__A1_N _16603_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24215_ _24214_/CLK _24215_/D HRESETn VGND VGND VPWR VPWR _24215_/Q sky130_fd_sc_hd__dfrtp_4
X_21427_ _21284_/A VGND VGND VPWR VPWR _21427_/X sky130_fd_sc_hd__buf_2
X_25195_ _23989_/CLK _14204_/X HRESETn VGND VGND VPWR VPWR _20506_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21739__B _21019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14922__A _14922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12160_ _25151_/Q _14338_/A _14339_/A _25152_/Q VGND VGND VPWR VPWR _12160_/X sky130_fd_sc_hd__and4_4
X_24146_ _24171_/CLK _18594_/X HRESETn VGND VGND VPWR VPWR _24146_/Q sky130_fd_sc_hd__dfrtp_4
X_21358_ _14212_/Y _14194_/A _14273_/Y _21548_/B VGND VGND VPWR VPWR _21359_/D sky130_fd_sc_hd__o22a_4
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23978__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_41_0_HCLK clkbuf_7_20_0_HCLK/X VGND VGND VPWR VPWR _23884_/CLK sky130_fd_sc_hd__clkbuf_1
X_20309_ _21801_/B _20304_/X _19988_/X _20304_/X VGND VGND VPWR VPWR _20309_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19057__B1 _19056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13538__A _25289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12091_ _12090_/Y _12086_/X _11867_/X _12073_/Y VGND VGND VPWR VPWR _12091_/X sky130_fd_sc_hd__a2bb2o_4
X_24077_ _24077_/CLK _24077_/D HRESETn VGND VGND VPWR VPWR _20427_/C sky130_fd_sc_hd__dfrtp_4
X_21289_ _16716_/A _21280_/B VGND VGND VPWR VPWR _21289_/X sky130_fd_sc_hd__or2_4
XFILLER_7_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21755__A _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23028_ _23027_/X VGND VGND VPWR VPWR _23028_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18804__B1 _18707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15618__B1 _11829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24941__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15850_ _15713_/A VGND VGND VPWR VPWR _15850_/X sky130_fd_sc_hd__buf_2
XFILLER_103_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14801_ _14815_/C _14801_/B _25037_/Q VGND VGND VPWR VPWR _14802_/B sky130_fd_sc_hd__or3_4
XFILLER_131_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15781_ _15728_/A VGND VGND VPWR VPWR _15781_/X sky130_fd_sc_hd__buf_2
X_12993_ _12993_/A _13107_/A _12292_/Y _12992_/Y VGND VGND VPWR VPWR _12993_/X sky130_fd_sc_hd__or4_4
XFILLER_45_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24979_ _24980_/CLK _24979_/D HRESETn VGND VGND VPWR VPWR _15083_/A sky130_fd_sc_hd__dfrtp_4
X_17520_ _25509_/Q _24280_/Q _11855_/Y _17662_/B VGND VGND VPWR VPWR _17520_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13273__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14732_ _25054_/Q _14707_/A _14731_/X VGND VGND VPWR VPWR _14732_/X sky130_fd_sc_hd__a21o_4
X_11944_ _11942_/Y _11935_/X _11943_/X _11935_/X VGND VGND VPWR VPWR _25493_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16043__B1 _11809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20914__B2 _20913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18783__B _18743_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17451_ _19219_/C VGND VGND VPWR VPWR _17451_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24766__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11875_ _11873_/X VGND VGND VPWR VPWR _11924_/A sky130_fd_sc_hd__inv_2
X_14663_ _19014_/B _19038_/C _19038_/D _14663_/D VGND VGND VPWR VPWR _14663_/X sky130_fd_sc_hd__and4_4
X_16402_ _15089_/Y _16400_/X _16401_/X _16400_/X VGND VGND VPWR VPWR _24588_/D sky130_fd_sc_hd__a2bb2o_4
X_13614_ _14641_/B _13613_/X _14641_/B _13613_/X VGND VGND VPWR VPWR _14792_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22667__A1 _16590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17382_ _17206_/X _17347_/B VGND VGND VPWR VPWR _17383_/C sky130_fd_sc_hd__nand2_4
X_14594_ _13576_/Y _14567_/B VGND VGND VPWR VPWR _14594_/Y sky130_fd_sc_hd__nand2_4
X_19121_ _19119_/Y _19120_/X _19077_/X _19120_/X VGND VGND VPWR VPWR _23839_/D sky130_fd_sc_hd__a2bb2o_4
X_16333_ _16332_/Y _16330_/X _16235_/X _16330_/X VGND VGND VPWR VPWR _24612_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13545_ _13543_/Y _13559_/A _22576_/A _25081_/Q VGND VGND VPWR VPWR _13554_/A sky130_fd_sc_hd__a2bb2o_4
X_19052_ _19052_/A VGND VGND VPWR VPWR _19052_/X sky130_fd_sc_hd__buf_2
XFILLER_51_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13476_ _13475_/X VGND VGND VPWR VPWR _13476_/Y sky130_fd_sc_hd__inv_2
X_16264_ _16263_/Y _16259_/X _15986_/X _16259_/X VGND VGND VPWR VPWR _24636_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18003_ _18010_/A VGND VGND VPWR VPWR _18046_/A sky130_fd_sc_hd__buf_2
X_12427_ _12410_/A _12424_/B _12427_/C VGND VGND VPWR VPWR _12427_/X sky130_fd_sc_hd__or3_4
X_15215_ _15065_/Y _15212_/X VGND VGND VPWR VPWR _15216_/C sky130_fd_sc_hd__or2_4
XFILLER_138_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15928__A _15674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19296__B1 _19294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16195_ _23232_/A VGND VGND VPWR VPWR _16195_/Y sky130_fd_sc_hd__inv_2
X_12358_ _25337_/Q VGND VGND VPWR VPWR _12358_/Y sky130_fd_sc_hd__inv_2
X_15146_ _15389_/A _24571_/Q _24991_/Q _15145_/Y VGND VGND VPWR VPWR _15146_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13448__A _13310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15077_ _15077_/A VGND VGND VPWR VPWR _15077_/Y sky130_fd_sc_hd__inv_2
X_19954_ _19954_/A VGND VGND VPWR VPWR _22245_/B sky130_fd_sc_hd__inv_2
XANTENNA__19048__B1 _18955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12289_ _12244_/Y _12252_/Y _12289_/C _12288_/X VGND VGND VPWR VPWR _12290_/B sky130_fd_sc_hd__or4_4
X_14028_ _13997_/X _13998_/X _14006_/A VGND VGND VPWR VPWR _14030_/A sky130_fd_sc_hd__o21ai_4
X_18905_ _22208_/B _18902_/X _16867_/X _18902_/X VGND VGND VPWR VPWR _18905_/X sky130_fd_sc_hd__a2bb2o_4
X_19885_ _19885_/A VGND VGND VPWR VPWR _19885_/X sky130_fd_sc_hd__buf_2
X_18836_ _16518_/A _24121_/Q _16518_/Y _18792_/B VGND VGND VPWR VPWR _18836_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15663__A _15670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18767_ _18767_/A _18767_/B VGND VGND VPWR VPWR _18767_/X sky130_fd_sc_hd__or2_4
X_15979_ _12204_/Y _15975_/X _15758_/X _15978_/X VGND VGND VPWR VPWR _24743_/D sky130_fd_sc_hd__a2bb2o_4
X_17718_ _17713_/X _21465_/A _17713_/X _21465_/A VGND VGND VPWR VPWR _18318_/B sky130_fd_sc_hd__a2bb2o_4
X_18698_ _18705_/A _18705_/B _18698_/C _18697_/X VGND VGND VPWR VPWR _18698_/X sky130_fd_sc_hd__or4_4
X_17649_ _17642_/A _17645_/B _17648_/X VGND VGND VPWR VPWR _17649_/X sky130_fd_sc_hd__and3_4
XFILLER_63_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13399__B2 _11964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24436__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20660_ _20659_/X VGND VGND VPWR VPWR _23981_/D sky130_fd_sc_hd__inv_2
X_19319_ _19317_/Y _19312_/X _19294_/X _19318_/X VGND VGND VPWR VPWR _23770_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22122__A3 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20591_ _25096_/Q _20443_/B VGND VGND VPWR VPWR _20591_/X sky130_fd_sc_hd__or2_4
XFILLER_31_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12527__A _12527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22330_ _21917_/X _22330_/B _22329_/X VGND VGND VPWR VPWR _22330_/X sky130_fd_sc_hd__and3_4
XFILLER_104_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20744__A _20761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22261_ _21260_/X _22241_/X _22256_/X _22259_/Y _22260_/X VGND VGND VPWR VPWR _22261_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__21559__B _13467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18214__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24000_ _24033_/CLK _24000_/D HRESETn VGND VGND VPWR VPWR _24000_/Q sky130_fd_sc_hd__dfrtp_4
X_21212_ _21015_/A VGND VGND VPWR VPWR _21220_/A sky130_fd_sc_hd__buf_2
XFILLER_133_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22192_ _22200_/A _22192_/B VGND VGND VPWR VPWR _22192_/X sky130_fd_sc_hd__or2_4
XANTENNA__15045__A2_N _24447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25295__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_0_0_HCLK clkbuf_8_1_0_HCLK/A VGND VGND VPWR VPWR _24398_/CLK sky130_fd_sc_hd__clkbuf_1
X_21143_ _21143_/A VGND VGND VPWR VPWR _21143_/X sky130_fd_sc_hd__buf_2
XFILLER_132_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16591__A1_N _16590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_28_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25224__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21575__A _16535_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21074_ _21005_/B _21074_/B VGND VGND VPWR VPWR _21074_/X sky130_fd_sc_hd__and2_4
XFILLER_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20025_ _22329_/B _20024_/X _19975_/X _20024_/X VGND VGND VPWR VPWR _20025_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23928__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24902_ _24487_/CLK _24902_/D HRESETn VGND VGND VPWR VPWR _15583_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_115_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11885__A1 _13678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21294__B _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24833_ _24868_/CLK _15804_/X HRESETn VGND VGND VPWR VPWR _24833_/Q sky130_fd_sc_hd__dfrtp_4
X_21976_ _18359_/Y _21977_/B _18348_/Y _20331_/A VGND VGND VPWR VPWR _21976_/X sky130_fd_sc_hd__o22a_4
X_24764_ _24792_/CLK _24764_/D HRESETn VGND VGND VPWR VPWR _24764_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16025__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20927_ _20925_/Y _20922_/Y _20931_/B VGND VGND VPWR VPWR _20927_/X sky130_fd_sc_hd__o21a_4
XPHY_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23715_ _23580_/CLK _19474_/X VGND VGND VPWR VPWR _23715_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24695_ _24699_/CLK _16099_/X HRESETn VGND VGND VPWR VPWR _23187_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17773__B1 _16955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ _11659_/Y _24225_/Q _11659_/Y _24225_/Q VGND VGND VPWR VPWR _11666_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20858_ _16697_/Y _20836_/X _20845_/X _20857_/X VGND VGND VPWR VPWR _20858_/X sky130_fd_sc_hd__o22a_4
XPHY_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23646_ _24186_/CLK _19679_/X VGND VGND VPWR VPWR _19678_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20806__A1_N _20680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23577_ _24926_/CLK _19876_/X VGND VGND VPWR VPWR _19875_/A sky130_fd_sc_hd__dfxtp_4
X_20789_ _20770_/X _20788_/X _24905_/Q _20774_/X VGND VGND VPWR VPWR _24022_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12243__A1_N _12430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _13395_/A _13330_/B VGND VGND VPWR VPWR _13330_/X sky130_fd_sc_hd__or2_4
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22528_ _15023_/A _22525_/X _22527_/X VGND VGND VPWR VPWR _22528_/X sky130_fd_sc_hd__o21a_4
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25316_ _25316_/CLK _25316_/D HRESETn VGND VGND VPWR VPWR _25316_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20654__A _25186_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _13440_/A _19067_/A VGND VGND VPWR VPWR _13261_/X sky130_fd_sc_hd__or2_4
XFILLER_127_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23030__A _23007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22459_ _22280_/X VGND VGND VPWR VPWR _22786_/A sky130_fd_sc_hd__buf_2
X_25247_ _25263_/CLK _25247_/D HRESETn VGND VGND VPWR VPWR _25247_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12212_ _12201_/X _12212_/B _12208_/X _12212_/D VGND VGND VPWR VPWR _12212_/X sky130_fd_sc_hd__or4_4
X_15000_ _15000_/A VGND VGND VPWR VPWR _15070_/B sky130_fd_sc_hd__buf_2
X_13192_ _13188_/X _13191_/X _13174_/X VGND VGND VPWR VPWR _13192_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12258__A1_N _12290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25178_ _25178_/CLK _25178_/D HRESETn VGND VGND VPWR VPWR _14261_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15839__B1 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12143_ _12143_/A VGND VGND VPWR VPWR _12143_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13268__A _13454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24129_ _24555_/CLK _24129_/D HRESETn VGND VGND VPWR VPWR _24129_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12074_ _12073_/Y VGND VGND VPWR VPWR _12074_/X sky130_fd_sc_hd__buf_2
X_16951_ _16946_/X _16947_/X _16949_/X _16950_/X VGND VGND VPWR VPWR _16952_/D sky130_fd_sc_hd__or4_4
XANTENNA__16579__A _24519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15902_ _12775_/Y _15900_/X _15620_/X _15900_/X VGND VGND VPWR VPWR _15902_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19670_ _19668_/Y _19663_/X _19645_/X _19669_/X VGND VGND VPWR VPWR _19670_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18497__C _18503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16882_ _16879_/Y _16880_/X _16881_/X _16880_/X VGND VGND VPWR VPWR _16882_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19450__B1 _19404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16264__B1 _15986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18621_ _24137_/Q VGND VGND VPWR VPWR _18675_/A sky130_fd_sc_hd__inv_2
X_15833_ _15829_/A VGND VGND VPWR VPWR _15833_/X sky130_fd_sc_hd__buf_2
XANTENNA__24947__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18552_ _18552_/A VGND VGND VPWR VPWR _18552_/Y sky130_fd_sc_hd__inv_2
X_15764_ _12563_/Y _15763_/X _15627_/X _15763_/X VGND VGND VPWR VPWR _24847_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12976_ _12976_/A _12979_/B VGND VGND VPWR VPWR _12977_/C sky130_fd_sc_hd__nand2_4
XANTENNA__16016__B1 _15949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17503_ _11776_/A _17630_/A _11756_/A _17600_/C VGND VGND VPWR VPWR _17505_/C sky130_fd_sc_hd__a2bb2o_4
X_14715_ _14714_/X VGND VGND VPWR VPWR _14716_/A sky130_fd_sc_hd__buf_2
X_11927_ _11923_/Y _11926_/X RsRx_S1 _11926_/X VGND VGND VPWR VPWR _11927_/X sky130_fd_sc_hd__a2bb2o_4
X_18483_ _24176_/Q _18483_/B VGND VGND VPWR VPWR _18485_/B sky130_fd_sc_hd__or2_4
X_15695_ _15694_/X VGND VGND VPWR VPWR _15695_/X sky130_fd_sc_hd__buf_2
XFILLER_2_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17434_ _24314_/Q VGND VGND VPWR VPWR _17434_/Y sky130_fd_sc_hd__inv_2
X_14646_ _18087_/A VGND VGND VPWR VPWR _14646_/X sky130_fd_sc_hd__buf_2
XFILLER_127_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11858_ _15986_/A VGND VGND VPWR VPWR _11858_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19505__B2 _19500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17365_ _17365_/A _17371_/A VGND VGND VPWR VPWR _17369_/B sky130_fd_sc_hd__or2_4
X_11789_ _11787_/Y _11785_/X _11788_/X _11785_/X VGND VGND VPWR VPWR _11789_/X sky130_fd_sc_hd__a2bb2o_4
X_14577_ _14558_/X _14579_/B _13568_/X _14586_/A VGND VGND VPWR VPWR _14577_/X sky130_fd_sc_hd__and4_4
XFILLER_14_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19104_ _13180_/B VGND VGND VPWR VPWR _19104_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16316_ _16288_/X VGND VGND VPWR VPWR _16316_/X sky130_fd_sc_hd__buf_2
X_13528_ _13514_/A _13526_/Y _13527_/X _13524_/B VGND VGND VPWR VPWR _13529_/A sky130_fd_sc_hd__a211o_4
X_17296_ _17239_/A _17293_/X VGND VGND VPWR VPWR _17296_/X sky130_fd_sc_hd__or2_4
X_19035_ _19034_/Y _19030_/X _19010_/X _19030_/A VGND VGND VPWR VPWR _19035_/X sky130_fd_sc_hd__a2bb2o_4
X_16247_ _16225_/A VGND VGND VPWR VPWR _16247_/X sky130_fd_sc_hd__buf_2
X_13459_ _13320_/A _13459_/B VGND VGND VPWR VPWR _13459_/X sky130_fd_sc_hd__or2_4
XFILLER_127_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16178_ _14772_/A _16176_/Y _13739_/B _16176_/Y VGND VGND VPWR VPWR _24666_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15129_ _15128_/Y _22608_/A _15128_/Y _22608_/A VGND VGND VPWR VPWR _15129_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19937_ _19935_/Y _19931_/X _19618_/X _19936_/X VGND VGND VPWR VPWR _19937_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19868_ _19880_/A VGND VGND VPWR VPWR _19868_/X sky130_fd_sc_hd__buf_2
XFILLER_110_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19441__B1 _19349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16255__B1 _16061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24688__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18819_ _18639_/Y _18783_/X VGND VGND VPWR VPWR _18819_/Y sky130_fd_sc_hd__nand2_4
X_19799_ _23605_/Q VGND VGND VPWR VPWR _21229_/B sky130_fd_sc_hd__inv_2
X_21830_ _21829_/Y _21143_/X _17427_/Y _17416_/A VGND VGND VPWR VPWR _21830_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24617__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21761_ _21616_/A _20158_/Y VGND VGND VPWR VPWR _21763_/B sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_4_3_0_HCLK_A clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18209__A _18177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21551__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20712_ _20712_/A VGND VGND VPWR VPWR _20713_/A sky130_fd_sc_hd__inv_2
XANTENNA__24270__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23500_ _23467_/CLK _23500_/D VGND VGND VPWR VPWR _20076_/A sky130_fd_sc_hd__dfxtp_4
X_24480_ _24496_/CLK _24480_/D HRESETn VGND VGND VPWR VPWR _24480_/Q sky130_fd_sc_hd__dfrtp_4
X_21692_ _21512_/X _21691_/X _21427_/X _25510_/Q _21428_/X VGND VGND VPWR VPWR _21692_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_52_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23431_ _23478_/CLK _20267_/X VGND VGND VPWR VPWR _20265_/A sky130_fd_sc_hd__dfxtp_4
X_20643_ _17396_/B _20643_/B _20651_/C VGND VGND VPWR VPWR _20643_/X sky130_fd_sc_hd__and3_4
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18648__A1_N _16565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21536__A1_N _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23362_ _21005_/X VGND VGND VPWR VPWR IRQ[8] sky130_fd_sc_hd__buf_2
X_20574_ _20574_/A _20571_/A VGND VGND VPWR VPWR _20575_/B sky130_fd_sc_hd__nand2_4
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22313_ _12106_/Y _12097_/X _18369_/Y _12071_/A VGND VGND VPWR VPWR _22313_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25476__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25101_ _25101_/CLK _14493_/X HRESETn VGND VGND VPWR VPWR _25101_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15568__A _15563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21289__B _21280_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23293_ _24532_/Q _22467_/X _22834_/X _23292_/X VGND VGND VPWR VPWR _23294_/C sky130_fd_sc_hd__a211o_4
XANTENNA__25405__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25032_ _25029_/CLK _25032_/D HRESETn VGND VGND VPWR VPWR _14813_/C sky130_fd_sc_hd__dfrtp_4
X_22244_ _21668_/A _22242_/X _22243_/X VGND VGND VPWR VPWR _22244_/X sky130_fd_sc_hd__and3_4
XFILLER_106_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22803__A1 _24550_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17783__A _17837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22175_ _14261_/Y _14257_/A _17420_/Y _17415_/A VGND VGND VPWR VPWR _22175_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16494__B1 _16408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21126_ _21350_/B _21125_/X _21116_/A VGND VGND VPWR VPWR _21126_/X sky130_fd_sc_hd__o21a_4
X_21057_ _21004_/B _21038_/B VGND VGND VPWR VPWR _21057_/X sky130_fd_sc_hd__and2_4
XFILLER_59_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19432__B1 _19407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23009__B _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_115_0_HCLK clkbuf_7_57_0_HCLK/X VGND VGND VPWR VPWR _24545_/CLK sky130_fd_sc_hd__clkbuf_1
X_20008_ _22014_/B _20002_/X _19981_/X _20007_/X VGND VGND VPWR VPWR _23530_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_178_0_HCLK clkbuf_7_89_0_HCLK/X VGND VGND VPWR VPWR _24290_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22319__B1 _20663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12830_ _12830_/A VGND VGND VPWR VPWR _12830_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24358__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24816_ _25330_/CLK _15828_/X HRESETn VGND VGND VPWR VPWR _24816_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12807__B1 _22660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12761_ _25355_/Q VGND VGND VPWR VPWR _12761_/Y sky130_fd_sc_hd__inv_2
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24747_ _24785_/CLK _24747_/D HRESETn VGND VGND VPWR VPWR _24747_/Q sky130_fd_sc_hd__dfrtp_4
X_21959_ _21962_/A _19597_/A _14613_/A _19601_/Y VGND VGND VPWR VPWR _21959_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13480__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _23952_/Q VGND VGND VPWR VPWR _14513_/A sky130_fd_sc_hd__inv_2
X_11712_ _15782_/B VGND VGND VPWR VPWR _15640_/B sky130_fd_sc_hd__inv_2
XANTENNA__17023__A _24632_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12664_/A VGND VGND VPWR VPWR _12698_/A sky130_fd_sc_hd__buf_2
X_15480_ _16720_/A VGND VGND VPWR VPWR _15480_/X sky130_fd_sc_hd__buf_2
XFILLER_43_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24678_ _24334_/CLK _24678_/D HRESETn VGND VGND VPWR VPWR _22556_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22864__A _22654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14430_/Y _14426_/X _14400_/X _14408_/Y VGND VGND VPWR VPWR _25125_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23629_ _23388_/CLK _23629_/D VGND VGND VPWR VPWR _19725_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22583__B _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ _16994_/A _17149_/Y VGND VGND VPWR VPWR _17150_/X sky130_fd_sc_hd__or2_4
XFILLER_122_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14362_ _25146_/Q _14351_/X _25145_/Q _14356_/X VGND VGND VPWR VPWR _14362_/X sky130_fd_sc_hd__o22a_4
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23993__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16101_ _16094_/A VGND VGND VPWR VPWR _16101_/X sky130_fd_sc_hd__buf_2
XFILLER_128_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _13450_/A _13313_/B _13313_/C VGND VGND VPWR VPWR _13313_/X sky130_fd_sc_hd__and3_4
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14293_ _13522_/D _14292_/Y _13643_/B VGND VGND VPWR VPWR _25169_/D sky130_fd_sc_hd__o21a_4
X_17081_ _17029_/A _17079_/X _17080_/Y VGND VGND VPWR VPWR _24385_/D sky130_fd_sc_hd__o21a_4
XANTENNA__21199__B _21333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23922__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21058__B1 _22664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12338__A2 _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25146__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13244_ _13390_/A _13244_/B _13243_/X VGND VGND VPWR VPWR _13244_/X sky130_fd_sc_hd__or3_4
X_16032_ _16031_/Y _16027_/X _15964_/X _16027_/X VGND VGND VPWR VPWR _16032_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18789__A _18789_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13175_ _13167_/X _13172_/X _13174_/X VGND VGND VPWR VPWR _13175_/X sky130_fd_sc_hd__o21a_4
XFILLER_112_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12126_ _24097_/Q _12126_/B VGND VGND VPWR VPWR _12127_/B sky130_fd_sc_hd__and2_4
X_17983_ _17982_/X _23739_/Q VGND VGND VPWR VPWR _17983_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_11_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_22_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__22558__B1 _25517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19722_ _19719_/Y _19720_/X _19721_/X _19720_/X VGND VGND VPWR VPWR _23631_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_74_0_HCLK clkbuf_7_75_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_74_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12057_ _12057_/A VGND VGND VPWR VPWR _19581_/B sky130_fd_sc_hd__inv_2
X_16934_ _16108_/Y _24268_/Q _16108_/Y _24268_/Q VGND VGND VPWR VPWR _16937_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15644__C _11731_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19653_ _19638_/Y VGND VGND VPWR VPWR _19653_/X sky130_fd_sc_hd__buf_2
XANTENNA__21943__A _21454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24781__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16865_ _20085_/A VGND VGND VPWR VPWR _16872_/A sky130_fd_sc_hd__buf_2
XFILLER_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18604_ _16560_/Y _18603_/X _16560_/Y _18603_/X VGND VGND VPWR VPWR _18605_/D sky130_fd_sc_hd__a2bb2o_4
X_15816_ _15728_/A VGND VGND VPWR VPWR _15816_/X sky130_fd_sc_hd__buf_2
XFILLER_24_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24099__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24710__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19584_ _21364_/C VGND VGND VPWR VPWR _19585_/A sky130_fd_sc_hd__buf_2
X_16796_ _16801_/A VGND VGND VPWR VPWR _16796_/X sky130_fd_sc_hd__buf_2
X_18535_ _18405_/Y _18539_/B _18534_/Y VGND VGND VPWR VPWR _18535_/X sky130_fd_sc_hd__o21a_4
XFILLER_80_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24028__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15747_ HWDATA[13] VGND VGND VPWR VPWR _15747_/X sky130_fd_sc_hd__buf_2
XFILLER_80_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12959_ _12959_/A _12959_/B VGND VGND VPWR VPWR _12960_/B sky130_fd_sc_hd__or2_4
XFILLER_34_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18466_ _18400_/Y _18524_/A _18523_/A VGND VGND VPWR VPWR _18466_/X sky130_fd_sc_hd__or3_4
X_15678_ _13540_/B VGND VGND VPWR VPWR _15684_/A sky130_fd_sc_hd__buf_2
X_17417_ _17432_/A VGND VGND VPWR VPWR _17417_/X sky130_fd_sc_hd__buf_2
XFILLER_33_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14629_ _14625_/Y _14628_/Y _14624_/X _14628_/A VGND VGND VPWR VPWR _25069_/D sky130_fd_sc_hd__o22a_4
X_18397_ _16223_/Y _18461_/A _16223_/Y _18461_/A VGND VGND VPWR VPWR _18404_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22493__B _22493_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17348_ _17348_/A _17348_/B VGND VGND VPWR VPWR _17371_/A sky130_fd_sc_hd__or2_4
XFILLER_14_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17279_ _17279_/A VGND VGND VPWR VPWR _17279_/X sky130_fd_sc_hd__buf_2
X_19018_ _19017_/X VGND VGND VPWR VPWR _19018_/X sky130_fd_sc_hd__buf_2
X_20290_ _20290_/A VGND VGND VPWR VPWR _20290_/X sky130_fd_sc_hd__buf_2
XANTENNA__22940__C _22812_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22261__A2 _22241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21837__B _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15818__A3 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24869__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23980_ _25219_/CLK _23980_/D HRESETn VGND VGND VPWR VPWR _23980_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21221__B1 _21211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22931_ _14927_/A _22929_/X _22524_/A _22930_/X VGND VGND VPWR VPWR _22932_/C sky130_fd_sc_hd__a211o_4
XFILLER_84_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24451__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22862_ _22861_/X VGND VGND VPWR VPWR _22862_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24601_ _24177_/CLK _24601_/D HRESETn VGND VGND VPWR VPWR _21531_/A sky130_fd_sc_hd__dfrtp_4
X_21813_ _21809_/X _21812_/X _21679_/X VGND VGND VPWR VPWR _21814_/C sky130_fd_sc_hd__o21a_4
XFILLER_71_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22793_ _13593_/X _21160_/X _22726_/B _22510_/A VGND VGND VPWR VPWR _22794_/A sky130_fd_sc_hd__a211o_4
XFILLER_58_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21744_ _21713_/Y _21744_/B _21737_/Y _21744_/D VGND VGND VPWR VPWR _21744_/X sky130_fd_sc_hd__or4_4
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24532_ _24561_/CLK _16548_/X HRESETn VGND VGND VPWR VPWR _24532_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22684__A _22425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17778__A _16916_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21675_ _21485_/A _21675_/B _21674_/X VGND VGND VPWR VPWR _21675_/X sky130_fd_sc_hd__and3_4
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24463_ _25016_/CLK _16732_/X HRESETn VGND VGND VPWR VPWR _24463_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20626_ _15465_/Y _20605_/X _20619_/X _20625_/X VGND VGND VPWR VPWR _20627_/A sky130_fd_sc_hd__a211o_4
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23414_ _23533_/CLK _20312_/X VGND VGND VPWR VPWR _20310_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_36_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24394_ _23478_/CLK _16886_/X HRESETn VGND VGND VPWR VPWR _20099_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23345_ _11970_/C _11967_/B _11959_/X VGND VGND VPWR VPWR _25540_/D sky130_fd_sc_hd__o21ai_4
X_20557_ _18874_/A _18874_/B VGND VGND VPWR VPWR _20557_/Y sky130_fd_sc_hd__nand2_4
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23276_ _23106_/X _23275_/X _21514_/X _24733_/Q _21520_/X VGND VGND VPWR VPWR _23276_/X
+ sky130_fd_sc_hd__a32o_4
X_20488_ _20488_/A _20488_/B VGND VGND VPWR VPWR _20488_/X sky130_fd_sc_hd__and2_4
X_22227_ _22009_/A _22227_/B VGND VGND VPWR VPWR _22227_/X sky130_fd_sc_hd__or2_4
X_25015_ _25024_/CLK _25015_/D HRESETn VGND VGND VPWR VPWR _25015_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_65_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22158_ _14386_/Y _21843_/X VGND VGND VPWR VPWR _22158_/Y sky130_fd_sc_hd__nor2_4
X_21109_ _24841_/Q _15649_/A _15655_/A _20674_/A _15658_/A VGND VGND VPWR VPWR _21109_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__19405__B1 _19404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23201__A1 _24561_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24539__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14980_ _25001_/Q VGND VGND VPWR VPWR _15267_/A sky130_fd_sc_hd__inv_2
X_22089_ _22089_/A _23082_/B VGND VGND VPWR VPWR _22093_/B sky130_fd_sc_hd__or2_4
XFILLER_93_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13931_ _13931_/A VGND VGND VPWR VPWR _13931_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16650_ _24494_/Q VGND VGND VPWR VPWR _16650_/Y sky130_fd_sc_hd__inv_2
X_13862_ _20466_/B VGND VGND VPWR VPWR _13862_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15601_ _15599_/Y _15600_/X _11800_/X _15600_/X VGND VGND VPWR VPWR _24895_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24121__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12813_ _12849_/A VGND VGND VPWR VPWR _12927_/A sky130_fd_sc_hd__buf_2
XFILLER_90_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16581_ _24518_/Q VGND VGND VPWR VPWR _16581_/Y sky130_fd_sc_hd__inv_2
X_13793_ _21996_/A VGND VGND VPWR VPWR _21498_/A sky130_fd_sc_hd__buf_2
XANTENNA__14377__A _15642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21515__A1 _21512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21515__B2 _21428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18320_ _18319_/X VGND VGND VPWR VPWR _18320_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13281__A _13156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15532_ _15531_/Y _15529_/X HADDR[6] _15529_/X VGND VGND VPWR VPWR _24918_/D sky130_fd_sc_hd__a2bb2o_4
X_12744_ _12859_/A VGND VGND VPWR VPWR _12744_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25398__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18251_ _11677_/Y _18249_/X _17424_/X _18249_/X VGND VGND VPWR VPWR _24218_/D sky130_fd_sc_hd__a2bb2o_4
X_15463_ _15476_/A VGND VGND VPWR VPWR _15463_/X sky130_fd_sc_hd__buf_2
XFILLER_128_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12675_ _12576_/Y _12674_/X VGND VGND VPWR VPWR _12689_/B sky130_fd_sc_hd__or2_4
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _17202_/A _17202_/B _17202_/C _17202_/D VGND VGND VPWR VPWR _17202_/X sky130_fd_sc_hd__or4_4
XANTENNA__25327__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ _15623_/A VGND VGND VPWR VPWR _14414_/X sky130_fd_sc_hd__buf_2
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18182_ _18150_/A _19348_/A VGND VGND VPWR VPWR _18182_/X sky130_fd_sc_hd__or2_4
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15394_ _15299_/A _15400_/B VGND VGND VPWR VPWR _15398_/B sky130_fd_sc_hd__or2_4
XFILLER_30_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ _17038_/B _17132_/X VGND VGND VPWR VPWR _17134_/B sky130_fd_sc_hd__or2_4
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ _14338_/Y _14344_/X VGND VGND VPWR VPWR _14345_/X sky130_fd_sc_hd__or2_4
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17064_ _17064_/A _17062_/X _17063_/X VGND VGND VPWR VPWR _17064_/X sky130_fd_sc_hd__and3_4
XANTENNA__21938__A _21458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14276_ _14275_/Y _14271_/X _13810_/X _14271_/A VGND VGND VPWR VPWR _25172_/D sky130_fd_sc_hd__a2bb2o_4
X_16015_ _16002_/X VGND VGND VPWR VPWR _16015_/X sky130_fd_sc_hd__buf_2
X_13227_ _13227_/A VGND VGND VPWR VPWR _13417_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12192__B1 _12290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24962__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13158_ _13186_/A _13158_/B VGND VGND VPWR VPWR _13158_/X sky130_fd_sc_hd__or2_4
XFILLER_97_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12109_ _25462_/Q VGND VGND VPWR VPWR _12109_/Y sky130_fd_sc_hd__inv_2
X_13089_ _12292_/Y _13087_/X _13088_/Y VGND VGND VPWR VPWR _13089_/X sky130_fd_sc_hd__o21a_4
X_17966_ _13610_/A VGND VGND VPWR VPWR _18024_/A sky130_fd_sc_hd__buf_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22769__A _22419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16917_ _16092_/A _16916_/A _16092_/Y _16916_/Y VGND VGND VPWR VPWR _16922_/B sky130_fd_sc_hd__o22a_4
X_19705_ _19683_/A _17472_/A _19219_/X VGND VGND VPWR VPWR _19705_/X sky130_fd_sc_hd__or3_4
XANTENNA__24209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17897_ _17904_/A _17896_/Y VGND VGND VPWR VPWR _17897_/X sky130_fd_sc_hd__and2_4
XANTENNA__16767__A _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22951__B1 _22090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16848_ _16801_/A VGND VGND VPWR VPWR _16848_/X sky130_fd_sc_hd__buf_2
X_19636_ _13159_/B VGND VGND VPWR VPWR _19636_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_161_0_HCLK clkbuf_7_80_0_HCLK/X VGND VGND VPWR VPWR _23683_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_4_0_HCLK clkbuf_6_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19567_ _19574_/A VGND VGND VPWR VPWR _19567_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_18_0_HCLK clkbuf_7_9_0_HCLK/X VGND VGND VPWR VPWR _25305_/CLK sky130_fd_sc_hd__clkbuf_1
X_16779_ _15028_/Y _16778_/X _16525_/X _16778_/X VGND VGND VPWR VPWR _16779_/X sky130_fd_sc_hd__a2bb2o_4
X_18518_ _18478_/X _18496_/X _18442_/Y VGND VGND VPWR VPWR _18518_/X sky130_fd_sc_hd__o21a_4
XFILLER_94_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19498_ _22249_/B _19495_/X _11934_/X _19495_/X VGND VGND VPWR VPWR _23707_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18449_ _18445_/X _18446_/X _18447_/X _18448_/X VGND VGND VPWR VPWR _18449_/X sky130_fd_sc_hd__or4_4
XFILLER_33_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25068__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21460_ _21460_/A _21460_/B _21460_/C VGND VGND VPWR VPWR _21460_/X sky130_fd_sc_hd__and3_4
XANTENNA__11758__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20411_ _13376_/B VGND VGND VPWR VPWR _20411_/Y sky130_fd_sc_hd__inv_2
X_21391_ _21391_/A _21389_/X _21390_/X VGND VGND VPWR VPWR _21391_/X sky130_fd_sc_hd__and3_4
XANTENNA__16007__A _24730_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23130_ _22798_/A VGND VGND VPWR VPWR _23130_/X sky130_fd_sc_hd__buf_2
X_20342_ _23402_/Q VGND VGND VPWR VPWR _20342_/Y sky130_fd_sc_hd__inv_2
X_23061_ _23133_/A _23058_/X _23061_/C VGND VGND VPWR VPWR _23066_/C sky130_fd_sc_hd__and3_4
X_20273_ _20272_/X VGND VGND VPWR VPWR _20273_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12183__B1 _12291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18222__A _18046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22012_ _22007_/X _22011_/X _21481_/X VGND VGND VPWR VPWR _22012_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_66_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21286__C _21290_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24632__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22679__A _22782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23963_ _24070_/CLK _20995_/X HRESETn VGND VGND VPWR VPWR _23963_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15581__A _15588_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22914_ _16673_/Y _22914_/B VGND VGND VPWR VPWR _22914_/X sky130_fd_sc_hd__and2_4
XFILLER_84_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23894_ _23905_/CLK _23894_/D VGND VGND VPWR VPWR _13409_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_99_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16621__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13813__B _13813_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22845_ _12792_/Y _21428_/X _22843_/X _12559_/Y _22844_/X VGND VGND VPWR VPWR _22845_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_72_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14197__A _20657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12789__A2 _24774_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22776_ _15791_/A _22774_/X _22485_/X _25523_/Q _22775_/X VGND VGND VPWR VPWR _22776_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_125_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25491__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24515_ _24517_/CLK _24515_/D HRESETn VGND VGND VPWR VPWR _16590_/A sky130_fd_sc_hd__dfrtp_4
X_21727_ _21727_/A VGND VGND VPWR VPWR _21727_/Y sky130_fd_sc_hd__inv_2
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25495_ _23394_/CLK _25495_/D HRESETn VGND VGND VPWR VPWR _11932_/A sky130_fd_sc_hd__dfrtp_4
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25420__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12460_ _12235_/X _12459_/X VGND VGND VPWR VPWR _12461_/A sky130_fd_sc_hd__or2_4
X_21658_ _21658_/A _19942_/Y VGND VGND VPWR VPWR _21659_/C sky130_fd_sc_hd__or2_4
X_24446_ _24462_/CLK _16766_/X HRESETn VGND VGND VPWR VPWR _24446_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12391_ _12391_/A _12391_/B VGND VGND VPWR VPWR _12391_/X sky130_fd_sc_hd__or2_4
X_20609_ _23969_/Q _17388_/B VGND VGND VPWR VPWR _20609_/Y sky130_fd_sc_hd__nand2_4
X_21589_ _21277_/Y VGND VGND VPWR VPWR _21589_/X sky130_fd_sc_hd__buf_2
XANTENNA__12445__A _12199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24377_ _24720_/CLK _24377_/D HRESETn VGND VGND VPWR VPWR _24377_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15537__A1_N _13496_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14130_ _14132_/A _14127_/X _14128_/Y _14129_/X VGND VGND VPWR VPWR _14130_/X sky130_fd_sc_hd__o22a_4
X_23328_ _24464_/Q _22654_/X _23172_/X VGND VGND VPWR VPWR _23328_/X sky130_fd_sc_hd__o21a_4
XFILLER_10_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20662__A _20662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14061_ _14006_/A _14057_/X _14060_/X VGND VGND VPWR VPWR _25229_/D sky130_fd_sc_hd__o21ai_4
XANTENNA__15756__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23259_ _23085_/A _23256_/X _23259_/C VGND VGND VPWR VPWR _23259_/X sky130_fd_sc_hd__and3_4
XANTENNA__12174__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13012_ _13012_/A _13023_/A _13002_/B _13001_/D VGND VGND VPWR VPWR _13013_/A sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_5_6_0_HCLK_A clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17820_ _16914_/Y _17824_/B _17819_/Y VGND VGND VPWR VPWR _17820_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17971__A _18087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24373__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16860__B1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25123__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17751_ _16911_/Y _17867_/A _17747_/X _17750_/X VGND VGND VPWR VPWR _17751_/X sky130_fd_sc_hd__or4_4
XANTENNA__21493__A _21821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24302__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14963_ _14954_/X _14963_/B _14963_/C _14962_/X VGND VGND VPWR VPWR _14984_/B sky130_fd_sc_hd__or4_4
XFILLER_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25186__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16702_ _24473_/Q VGND VGND VPWR VPWR _16702_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15491__A _15490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13914_ _13895_/X _13927_/D _13909_/X _13892_/A VGND VGND VPWR VPWR _13914_/X sky130_fd_sc_hd__or4_4
X_17682_ _17665_/X _17682_/B _17681_/X VGND VGND VPWR VPWR _17682_/X sky130_fd_sc_hd__and3_4
X_14894_ _14893_/Y VGND VGND VPWR VPWR _15197_/A sky130_fd_sc_hd__buf_2
XFILLER_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19421_ _19419_/Y _19415_/X _19420_/X _19401_/A VGND VGND VPWR VPWR _19421_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16612__B1 _16528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16633_ _13741_/C _16632_/Y _16627_/X VGND VGND VPWR VPWR _24500_/D sky130_fd_sc_hd__o21a_4
XFILLER_62_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_234_0_HCLK clkbuf_8_235_0_HCLK/A VGND VGND VPWR VPWR _25368_/CLK sky130_fd_sc_hd__clkbuf_1
X_13845_ _13565_/Y _13843_/X _13803_/X _13843_/X VGND VGND VPWR VPWR _25244_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25508__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19352_ _19351_/Y _19346_/X _19307_/X _19333_/Y VGND VGND VPWR VPWR _19352_/X sky130_fd_sc_hd__a2bb2o_4
X_16564_ _16562_/Y _16558_/X _16393_/X _16563_/X VGND VGND VPWR VPWR _16564_/X sky130_fd_sc_hd__a2bb2o_4
X_13776_ _13775_/X VGND VGND VPWR VPWR _13784_/C sky130_fd_sc_hd__buf_2
XANTENNA__11819__A1_N _11815_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18303_ _21465_/A _18303_/B VGND VGND VPWR VPWR _18303_/X sky130_fd_sc_hd__and2_4
X_15515_ _11728_/B VGND VGND VPWR VPWR _15515_/Y sky130_fd_sc_hd__inv_2
X_12727_ _12726_/X VGND VGND VPWR VPWR _25392_/D sky130_fd_sc_hd__inv_2
X_19283_ _21235_/B _19278_/X _18919_/X _19278_/A VGND VGND VPWR VPWR _19283_/X sky130_fd_sc_hd__a2bb2o_4
X_16495_ _24551_/Q VGND VGND VPWR VPWR _16495_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18234_ _11664_/Y _18233_/X _15743_/X _18233_/X VGND VGND VPWR VPWR _18234_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15446_ _15446_/A VGND VGND VPWR VPWR _15446_/X sky130_fd_sc_hd__buf_2
X_12658_ _12651_/B VGND VGND VPWR VPWR _12659_/B sky130_fd_sc_hd__inv_2
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18165_ _18133_/A _18165_/B VGND VGND VPWR VPWR _18165_/X sky130_fd_sc_hd__or2_4
XFILLER_102_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15377_ _15376_/X VGND VGND VPWR VPWR _24977_/D sky130_fd_sc_hd__inv_2
XFILLER_8_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12589_ _12580_/X _12583_/X _12589_/C _12588_/X VGND VGND VPWR VPWR _12599_/C sky130_fd_sc_hd__or4_4
XFILLER_11_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22771__B _22626_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17116_ _17033_/D _17091_/X _17067_/X _17114_/B VGND VGND VPWR VPWR _17116_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16679__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14328_ _25156_/Q _12163_/X _14327_/Y VGND VGND VPWR VPWR _14328_/X sky130_fd_sc_hd__o21a_4
X_18096_ _18058_/A _18096_/B _18095_/X VGND VGND VPWR VPWR _18096_/X sky130_fd_sc_hd__or3_4
XFILLER_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17047_ _17047_/A _17091_/B VGND VGND VPWR VPWR _17048_/D sky130_fd_sc_hd__or2_4
XANTENNA__15666__A _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14259_ _14271_/A VGND VGND VPWR VPWR _14259_/X sky130_fd_sc_hd__buf_2
XFILLER_125_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24325__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18977__A _16786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18998_ _18988_/Y VGND VGND VPWR VPWR _18998_/X sky130_fd_sc_hd__buf_2
XFILLER_100_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16851__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24043__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_44_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_44_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17949_ _17930_/A _20209_/A VGND VGND VPWR VPWR _17950_/C sky130_fd_sc_hd__or2_4
XANTENNA__16497__A _24550_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22924__B1 _22798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20960_ _12125_/A _12163_/B VGND VGND VPWR VPWR _24095_/D sky130_fd_sc_hd__nor2_4
XFILLER_61_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19619_ _19628_/A VGND VGND VPWR VPWR _19619_/X sky130_fd_sc_hd__buf_2
X_20891_ _20882_/X _20890_/X _24482_/Q _20886_/X VGND VGND VPWR VPWR _20891_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25249__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21850__B _21220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22630_ _21064_/A _22627_/X _21098_/X _22629_/X VGND VGND VPWR VPWR _22630_/Y sky130_fd_sc_hd__a22oi_4
X_22561_ _21105_/A _22559_/X _22103_/X _22560_/X VGND VGND VPWR VPWR _22562_/B sky130_fd_sc_hd__o22a_4
XANTENNA__14745__A _14744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18217__A _18217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21512_ _21511_/X VGND VGND VPWR VPWR _21512_/X sky130_fd_sc_hd__buf_2
XFILLER_33_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24300_ _25436_/CLK _17623_/Y HRESETn VGND VGND VPWR VPWR _17543_/A sky130_fd_sc_hd__dfrtp_4
X_22492_ _22490_/X _22492_/B _22440_/C VGND VGND VPWR VPWR _22492_/X sky130_fd_sc_hd__or3_4
X_25280_ _24252_/CLK _13706_/X HRESETn VGND VGND VPWR VPWR _13693_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_72_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21443_ _22792_/A _21421_/Y _21436_/Y _21437_/X _21442_/X VGND VGND VPWR VPWR _21444_/A
+ sky130_fd_sc_hd__a32o_4
X_24231_ _23826_/CLK _24231_/D HRESETn VGND VGND VPWR VPWR _24231_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21578__A _15668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24162_ _24162_/CLK _24162_/D HRESETn VGND VGND VPWR VPWR _24162_/Q sky130_fd_sc_hd__dfrtp_4
X_21374_ _14691_/A _21374_/B _21374_/C VGND VGND VPWR VPWR _21374_/X sky130_fd_sc_hd__and3_4
XANTENNA__24884__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20325_ _23408_/Q VGND VGND VPWR VPWR _21968_/A sky130_fd_sc_hd__inv_2
X_23113_ _23105_/X _23109_/Y _22863_/X _23112_/X VGND VGND VPWR VPWR _23113_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24813__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24093_ _25309_/CLK MSI_S2 HRESETn VGND VGND VPWR VPWR _24093_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12156__B1 _12092_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_126_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_126_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23044_ _21416_/A VGND VGND VPWR VPWR _23044_/X sky130_fd_sc_hd__buf_2
X_20256_ _23435_/Q VGND VGND VPWR VPWR _22189_/B sky130_fd_sc_hd__inv_2
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20187_ _20186_/Y _20182_/X _20123_/X _20182_/A VGND VGND VPWR VPWR _20187_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16842__B1 _16604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21744__C _21737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24995_ _24995_/CLK _15288_/X HRESETn VGND VGND VPWR VPWR _24995_/Q sky130_fd_sc_hd__dfrtp_4
X_11960_ _17445_/C VGND VGND VPWR VPWR _11967_/B sky130_fd_sc_hd__inv_2
XFILLER_131_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23946_ _25199_/CLK _23945_/Q HRESETn VGND VGND VPWR VPWR _23946_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11891_ _11869_/B VGND VGND VPWR VPWR _11892_/A sky130_fd_sc_hd__inv_2
X_23877_ _23869_/CLK _23877_/D VGND VGND VPWR VPWR _19009_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13630_ _13630_/A VGND VGND VPWR VPWR _17928_/A sky130_fd_sc_hd__buf_2
X_22828_ _16678_/Y _22790_/A _15595_/Y _22827_/X VGND VGND VPWR VPWR _22828_/X sky130_fd_sc_hd__o22a_4
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20657__A _20657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_64_0_HCLK clkbuf_8_65_0_HCLK/A VGND VGND VPWR VPWR _25098_/CLK sky130_fd_sc_hd__clkbuf_1
X_13561_ _25247_/Q _13559_/Y _13544_/A _14572_/A VGND VGND VPWR VPWR _13564_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22759_ _21108_/B VGND VGND VPWR VPWR _22759_/X sky130_fd_sc_hd__buf_2
X_15300_ _24973_/Q VGND VGND VPWR VPWR _15301_/D sky130_fd_sc_hd__inv_2
X_12512_ _25419_/Q VGND VGND VPWR VPWR _12512_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16280_ _16280_/A VGND VGND VPWR VPWR _16280_/X sky130_fd_sc_hd__buf_2
XFILLER_38_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13492_ _13491_/Y _13489_/X _11862_/X _13489_/X VGND VGND VPWR VPWR _25305_/D sky130_fd_sc_hd__a2bb2o_4
X_25478_ _25478_/CLK _25478_/D HRESETn VGND VGND VPWR VPWR _25478_/Q sky130_fd_sc_hd__dfrtp_4
X_15231_ _15210_/B _15210_/C VGND VGND VPWR VPWR _15232_/A sky130_fd_sc_hd__or2_4
XFILLER_90_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12443_ _12440_/C _12432_/B VGND VGND VPWR VPWR _12447_/A sky130_fd_sc_hd__or2_4
XANTENNA__17966__A _13610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24429_ _24431_/CLK _24429_/D HRESETn VGND VGND VPWR VPWR _24429_/Q sky130_fd_sc_hd__dfrtp_4
X_15162_ _15132_/X _15162_/B _15162_/C _15161_/X VGND VGND VPWR VPWR _15162_/X sky130_fd_sc_hd__or4_4
X_12374_ _12374_/A VGND VGND VPWR VPWR _12374_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14113_ _23950_/Q _14098_/X _14099_/A VGND VGND VPWR VPWR _14113_/X sky130_fd_sc_hd__or3_4
XFILLER_125_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24554__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15093_ _15092_/Y _16445_/A _15092_/Y _16445_/A VGND VGND VPWR VPWR _15093_/X sky130_fd_sc_hd__a2bb2o_4
X_19970_ _19970_/A VGND VGND VPWR VPWR _22348_/B sky130_fd_sc_hd__inv_2
XFILLER_125_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12903__A _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14044_ _13982_/A _13983_/X _13984_/A _13980_/A VGND VGND VPWR VPWR _14045_/B sky130_fd_sc_hd__or4_4
X_18921_ _23908_/Q VGND VGND VPWR VPWR _18921_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13718__B _13686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18797__A _18630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18852_ _16520_/Y _18623_/A _16520_/Y _18623_/A VGND VGND VPWR VPWR _18852_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16833__B1 _15747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17803_ _17738_/X _17794_/B _17802_/X VGND VGND VPWR VPWR _17803_/X sky130_fd_sc_hd__and3_4
X_18783_ _18680_/D _18743_/C VGND VGND VPWR VPWR _18783_/X sky130_fd_sc_hd__or2_4
XFILLER_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15995_ _15995_/A VGND VGND VPWR VPWR _15995_/X sky130_fd_sc_hd__buf_2
X_17734_ _17734_/A VGND VGND VPWR VPWR _17734_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12060__D _12059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14946_ _14990_/A _14944_/Y _25000_/Q _14945_/Y VGND VGND VPWR VPWR _14946_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15652__C _11732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17665_ _17494_/Y _17685_/A VGND VGND VPWR VPWR _17665_/X sky130_fd_sc_hd__or2_4
X_14877_ _14798_/B _14872_/B _14872_/Y VGND VGND VPWR VPWR _14877_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22119__D1 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25342__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16616_ _16616_/A VGND VGND VPWR VPWR _16616_/Y sky130_fd_sc_hd__inv_2
X_19404_ _19642_/A VGND VGND VPWR VPWR _19404_/X sky130_fd_sc_hd__buf_2
X_13828_ _22576_/A _13825_/X _11818_/X _13825_/X VGND VGND VPWR VPWR _25253_/D sky130_fd_sc_hd__a2bb2o_4
X_17596_ _17515_/A _17596_/B VGND VGND VPWR VPWR _17596_/X sky130_fd_sc_hd__or2_4
X_16547_ _24532_/Q VGND VGND VPWR VPWR _16547_/Y sky130_fd_sc_hd__inv_2
X_19335_ _19331_/Y _19334_/X _19313_/X _19334_/X VGND VGND VPWR VPWR _23764_/D sky130_fd_sc_hd__a2bb2o_4
X_13759_ _13759_/A VGND VGND VPWR VPWR _13759_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20145__B1 _20123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19266_ _19278_/A VGND VGND VPWR VPWR _19266_/X sky130_fd_sc_hd__buf_2
X_16478_ _24558_/Q VGND VGND VPWR VPWR _16478_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22782__A _22782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18217_ _18217_/A _18217_/B _18217_/C VGND VGND VPWR VPWR _18217_/X sky130_fd_sc_hd__or3_4
X_15429_ _13950_/X _15429_/B _13963_/X _14245_/X VGND VGND VPWR VPWR _15435_/A sky130_fd_sc_hd__or4_4
X_19197_ _19197_/A VGND VGND VPWR VPWR _19197_/X sky130_fd_sc_hd__buf_2
XFILLER_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18148_ _18180_/A _23863_/Q VGND VGND VPWR VPWR _18149_/C sky130_fd_sc_hd__or2_4
XFILLER_8_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24295__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18079_ _18079_/A VGND VGND VPWR VPWR _18097_/A sky130_fd_sc_hd__buf_2
XFILLER_105_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20110_ _20110_/A VGND VGND VPWR VPWR _20110_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24224__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21090_ _21729_/A _21089_/Y _24631_/Q _21729_/A VGND VGND VPWR VPWR _21090_/X sky130_fd_sc_hd__a2bb2o_4
X_20041_ _20040_/Y _20036_/X _20019_/X _20036_/A VGND VGND VPWR VPWR _20041_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23118__A _22782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23800_ _23798_/CLK _19233_/X VGND VGND VPWR VPWR _13340_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24083__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24780_ _24780_/CLK _15901_/X HRESETn VGND VGND VPWR VPWR _24780_/Q sky130_fd_sc_hd__dfrtp_4
X_21992_ _21989_/Y _21990_/X _21978_/X _21991_/X VGND VGND VPWR VPWR _23340_/B sky130_fd_sc_hd__a211o_4
XANTENNA__21861__A _23085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12348__A2_N _24819_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23731_ _23887_/CLK _23731_/D VGND VGND VPWR VPWR _17985_/B sky130_fd_sc_hd__dfxtp_4
X_20943_ _20943_/A _24057_/Q _13666_/X VGND VGND VPWR VPWR _20943_/X sky130_fd_sc_hd__or3_4
XPHY_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22676__B _22913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25083__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ _23398_/CLK _19633_/X VGND VGND VPWR VPWR _19631_/A sky130_fd_sc_hd__dfxtp_4
X_20874_ _13663_/A _13663_/B VGND VGND VPWR VPWR _20879_/B sky130_fd_sc_hd__or2_4
XPHY_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25012__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25401_ _25400_/CLK _25401_/D HRESETn VGND VGND VPWR VPWR _12570_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22613_ _24225_/Q _22613_/B VGND VGND VPWR VPWR _22613_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__20136__B1 _20089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14475__A _21027_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23593_ _23581_/CLK _19832_/X VGND VGND VPWR VPWR _23593_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17001__B1 _24724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25332_ _25351_/CLK _13091_/X HRESETn VGND VGND VPWR VPWR _12992_/A sky130_fd_sc_hd__dfrtp_4
X_22544_ _22123_/A VGND VGND VPWR VPWR _22544_/X sky130_fd_sc_hd__buf_2
XANTENNA__23086__C1 _23085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25263_ _25263_/CLK _13785_/X HRESETn VGND VGND VPWR VPWR _25263_/Q sky130_fd_sc_hd__dfrtp_4
X_22475_ _22419_/X VGND VGND VPWR VPWR _22475_/X sky130_fd_sc_hd__buf_2
XFILLER_6_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24214_ _24214_/CLK _18257_/X HRESETn VGND VGND VPWR VPWR _24214_/Q sky130_fd_sc_hd__dfrtp_4
X_21426_ _21426_/A _22998_/A VGND VGND VPWR VPWR _21426_/X sky130_fd_sc_hd__or2_4
XFILLER_136_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25194_ _23989_/CLK _14206_/X HRESETn VGND VGND VPWR VPWR _14205_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17503__A1_N _11776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21357_ _21139_/B VGND VGND VPWR VPWR _21548_/B sky130_fd_sc_hd__buf_2
X_24145_ _24171_/CLK _18596_/Y HRESETn VGND VGND VPWR VPWR _24145_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20308_ _20308_/A VGND VGND VPWR VPWR _21801_/B sky130_fd_sc_hd__inv_2
XFILLER_122_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12090_ _12090_/A VGND VGND VPWR VPWR _12090_/Y sky130_fd_sc_hd__inv_2
X_21288_ _21287_/Y VGND VGND VPWR VPWR _21302_/A sky130_fd_sc_hd__buf_2
XFILLER_104_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24076_ _25137_/CLK _24076_/D HRESETn VGND VGND VPWR VPWR _20445_/B sky130_fd_sc_hd__dfstp_4
X_20239_ _20237_/Y _20233_/X _19758_/X _20238_/X VGND VGND VPWR VPWR _23442_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23027_ _22753_/X _23025_/X _22684_/X _23026_/X VGND VGND VPWR VPWR _23027_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16815__B1 HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23947__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14800_ _14814_/C _14799_/X _25035_/Q VGND VGND VPWR VPWR _14801_/B sky130_fd_sc_hd__or3_4
X_15780_ _15552_/Y _15669_/X _15774_/X _24839_/Q _15779_/X VGND VGND VPWR VPWR _15780_/X
+ sky130_fd_sc_hd__a32o_4
X_12992_ _12992_/A VGND VGND VPWR VPWR _12992_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24978_ _24980_/CLK _24978_/D HRESETn VGND VGND VPWR VPWR _15374_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14731_ _14726_/X _14730_/Y _14723_/Y VGND VGND VPWR VPWR _14731_/X sky130_fd_sc_hd__a21o_4
X_11943_ _19622_/A VGND VGND VPWR VPWR _11943_/X sky130_fd_sc_hd__buf_2
X_23929_ _25098_/CLK _20977_/B HRESETn VGND VGND VPWR VPWR _14096_/C sky130_fd_sc_hd__dfstp_4
XFILLER_72_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17450_ _17449_/X VGND VGND VPWR VPWR _19219_/C sky130_fd_sc_hd__buf_2
XFILLER_44_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14662_ _25061_/Q VGND VGND VPWR VPWR _14663_/D sky130_fd_sc_hd__buf_2
XFILLER_17_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11874_ _25506_/Q _11869_/X _11873_/X VGND VGND VPWR VPWR _11874_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_33_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16401_ HWDATA[21] VGND VGND VPWR VPWR _16401_/X sky130_fd_sc_hd__buf_2
X_13613_ _25058_/Q VGND VGND VPWR VPWR _13613_/X sky130_fd_sc_hd__buf_2
X_17381_ _17370_/A _17381_/B _17380_/Y VGND VGND VPWR VPWR _24330_/D sky130_fd_sc_hd__and3_4
X_14593_ _14569_/A _14586_/X _14592_/Y _14590_/X _25079_/Q VGND VGND VPWR VPWR _14593_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22667__A2 _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13801__B1 _13800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19120_ _19106_/Y VGND VGND VPWR VPWR _19120_/X sky130_fd_sc_hd__buf_2
XFILLER_41_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16332_ _24612_/Q VGND VGND VPWR VPWR _16332_/Y sky130_fd_sc_hd__inv_2
X_13544_ _13544_/A VGND VGND VPWR VPWR _22576_/A sky130_fd_sc_hd__inv_2
X_19051_ _23863_/Q VGND VGND VPWR VPWR _19051_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16263_ _24636_/Q VGND VGND VPWR VPWR _16263_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24735__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13475_ _12066_/X _12072_/D _13533_/A _13533_/B VGND VGND VPWR VPWR _13475_/X sky130_fd_sc_hd__or4_4
Xclkbuf_6_8_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18002_ _18221_/A _18002_/B VGND VGND VPWR VPWR _18002_/X sky130_fd_sc_hd__or2_4
X_15214_ _14903_/X _15214_/B VGND VGND VPWR VPWR _15216_/B sky130_fd_sc_hd__or2_4
X_12426_ _12288_/X _12391_/B _12252_/Y VGND VGND VPWR VPWR _12427_/C sky130_fd_sc_hd__o21a_4
X_16194_ _16191_/Y _16187_/X _15940_/X _16193_/X VGND VGND VPWR VPWR _24663_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15145_ _24595_/Q VGND VGND VPWR VPWR _15145_/Y sky130_fd_sc_hd__inv_2
X_12357_ _13061_/A _24824_/Q _25343_/Q _12308_/Y VGND VGND VPWR VPWR _12360_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15076_ _15313_/A _24598_/Q _15313_/A _24598_/Q VGND VGND VPWR VPWR _15082_/B sky130_fd_sc_hd__a2bb2o_4
X_19953_ _19949_/Y _19952_/X _19612_/X _19952_/X VGND VGND VPWR VPWR _23548_/D sky130_fd_sc_hd__a2bb2o_4
X_12288_ _12283_/X _12287_/X VGND VGND VPWR VPWR _12288_/X sky130_fd_sc_hd__or2_4
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14027_ _13995_/B _14021_/X _14026_/Y VGND VGND VPWR VPWR _14070_/A sky130_fd_sc_hd__a21o_4
X_18904_ _23915_/Q VGND VGND VPWR VPWR _22208_/B sky130_fd_sc_hd__inv_2
XANTENNA__15944__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19884_ _19884_/A VGND VGND VPWR VPWR _21184_/B sky130_fd_sc_hd__inv_2
XFILLER_67_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18835_ _24563_/Q _24142_/Q _16465_/Y _18705_/A VGND VGND VPWR VPWR _18838_/B sky130_fd_sc_hd__o22a_4
XFILLER_68_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25523__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15978_ _15937_/Y VGND VGND VPWR VPWR _15978_/X sky130_fd_sc_hd__buf_2
X_18766_ _18765_/X VGND VGND VPWR VPWR _18767_/B sky130_fd_sc_hd__inv_2
XANTENNA__21158__A2 _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21681__A _21681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14929_ _15179_/A VGND VGND VPWR VPWR _15180_/A sky130_fd_sc_hd__inv_2
X_17717_ _17717_/A VGND VGND VPWR VPWR _21465_/A sky130_fd_sc_hd__buf_2
XFILLER_58_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18697_ _18743_/C _18704_/A VGND VGND VPWR VPWR _18697_/X sky130_fd_sc_hd__or2_4
XFILLER_63_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17648_ _17565_/A _17648_/B VGND VGND VPWR VPWR _17648_/X sky130_fd_sc_hd__or2_4
X_17579_ _17572_/X _17575_/X _17579_/C VGND VGND VPWR VPWR _17653_/B sky130_fd_sc_hd__or3_4
XFILLER_17_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12808__A _12896_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20669__A1 _20663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19318_ _19311_/Y VGND VGND VPWR VPWR _19318_/X sky130_fd_sc_hd__buf_2
X_20590_ _14452_/X _20589_/X VGND VGND VPWR VPWR _23944_/D sky130_fd_sc_hd__nor2_4
XFILLER_17_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24476__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19249_ _19256_/A VGND VGND VPWR VPWR _19249_/X sky130_fd_sc_hd__buf_2
X_22260_ _11661_/Y _21495_/X _21502_/A VGND VGND VPWR VPWR _22260_/X sky130_fd_sc_hd__a21o_4
XFILLER_118_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24405__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21211_ _22790_/A VGND VGND VPWR VPWR _21211_/X sky130_fd_sc_hd__buf_2
XANTENNA__21094__A1 _16075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17298__B1 _17279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22191_ _22078_/X _22189_/X _22191_/C VGND VGND VPWR VPWR _22191_/X sky130_fd_sc_hd__and3_4
X_21142_ _21142_/A VGND VGND VPWR VPWR _21142_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18863__A1_N _24560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21073_ _24735_/Q _21073_/B VGND VGND VPWR VPWR _21073_/X sky130_fd_sc_hd__or2_4
XANTENNA__15854__A _22835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21575__B _22695_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20024_ _20036_/A VGND VGND VPWR VPWR _20024_/X sky130_fd_sc_hd__buf_2
XFILLER_86_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22594__B2 _22593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24901_ _24487_/CLK _24901_/D HRESETn VGND VGND VPWR VPWR _24901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25264__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24832_ _24832_/CLK _15805_/X HRESETn VGND VGND VPWR VPWR _24832_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_14_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_55_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24763_ _25374_/CLK _15943_/X HRESETn VGND VGND VPWR VPWR _23210_/A sky130_fd_sc_hd__dfrtp_4
X_21975_ _21972_/X _21973_/X _21974_/X VGND VGND VPWR VPWR _21975_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__12834__B2 _24775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23714_ _23714_/CLK _23714_/D VGND VGND VPWR VPWR _19475_/A sky130_fd_sc_hd__dfxtp_4
X_20926_ _24054_/Q _24053_/Q _20922_/B VGND VGND VPWR VPWR _20931_/B sky130_fd_sc_hd__or3_4
XPHY_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24694_ _25354_/CLK _16102_/X HRESETn VGND VGND VPWR VPWR _24694_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18970__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23645_ _24186_/CLK _19681_/X VGND VGND VPWR VPWR _23645_/Q sky130_fd_sc_hd__dfxtp_4
X_20857_ _20856_/Y _20852_/X _13659_/X VGND VGND VPWR VPWR _20857_/X sky130_fd_sc_hd__o21a_4
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23576_ _23711_/CLK _19878_/X VGND VGND VPWR VPWR _23576_/Q sky130_fd_sc_hd__dfxtp_4
X_20788_ _20786_/Y _20783_/Y _20787_/X VGND VGND VPWR VPWR _20788_/X sky130_fd_sc_hd__o21a_4
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21704__A1_N _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25315_ _23377_/CLK _25315_/D HRESETn VGND VGND VPWR VPWR _25315_/Q sky130_fd_sc_hd__dfrtp_4
X_22527_ _22526_/X VGND VGND VPWR VPWR _22527_/X sky130_fd_sc_hd__buf_2
XANTENNA__15536__B1 HADDR[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20654__B _17404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_138_0_HCLK clkbuf_7_69_0_HCLK/X VGND VGND VPWR VPWR _25503_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13260_ _24191_/Q VGND VGND VPWR VPWR _13260_/X sky130_fd_sc_hd__buf_2
XANTENNA__23030__B _23030_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24146__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25246_ _25246_/CLK _13842_/X HRESETn VGND VGND VPWR VPWR _21952_/A sky130_fd_sc_hd__dfrtp_4
X_22458_ _22783_/A _22458_/B VGND VGND VPWR VPWR _22462_/C sky130_fd_sc_hd__nor2_4
XFILLER_109_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23074__A2 _21021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12211_ _25427_/Q _22400_/A _12209_/Y _12210_/Y VGND VGND VPWR VPWR _12212_/D sky130_fd_sc_hd__o22a_4
X_21409_ _21409_/A VGND VGND VPWR VPWR _22792_/A sky130_fd_sc_hd__buf_2
XANTENNA__22282__B1 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13191_ _13191_/A _13189_/X _13190_/X VGND VGND VPWR VPWR _13191_/X sky130_fd_sc_hd__and3_4
X_25177_ _23959_/CLK _25177_/D HRESETn VGND VGND VPWR VPWR _14263_/A sky130_fd_sc_hd__dfrtp_4
X_22389_ _22389_/A _22389_/B VGND VGND VPWR VPWR _22389_/X sky130_fd_sc_hd__or2_4
XFILLER_136_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12142_ _12127_/A _12127_/B _12141_/Y VGND VGND VPWR VPWR _12143_/A sky130_fd_sc_hd__o21a_4
X_24128_ _24133_/CLK _24128_/D HRESETn VGND VGND VPWR VPWR _24128_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12073_ _12072_/X VGND VGND VPWR VPWR _12073_/Y sky130_fd_sc_hd__inv_2
X_16950_ _16151_/Y _22181_/A _16159_/Y _24248_/Q VGND VGND VPWR VPWR _16950_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24059_ _24492_/CLK _24059_/D HRESETn VGND VGND VPWR VPWR _13667_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_42_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15901_ _12769_/Y _15896_/X _15758_/X _15900_/X VGND VGND VPWR VPWR _15901_/X sky130_fd_sc_hd__a2bb2o_4
X_16881_ _19790_/A VGND VGND VPWR VPWR _16881_/X sky130_fd_sc_hd__buf_2
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15832_ _12296_/Y _15829_/X _15623_/X _15829_/X VGND VGND VPWR VPWR _24813_/D sky130_fd_sc_hd__a2bb2o_4
X_18620_ _16603_/A _24121_/Q _16603_/Y _18619_/Y VGND VGND VPWR VPWR _18620_/X sky130_fd_sc_hd__o22a_4
XFILLER_77_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15763_ _15763_/A VGND VGND VPWR VPWR _15763_/X sky130_fd_sc_hd__buf_2
X_18551_ _18468_/Y _18550_/X VGND VGND VPWR VPWR _18552_/A sky130_fd_sc_hd__or2_4
X_12975_ _12964_/A _12975_/B _12974_/Y VGND VGND VPWR VPWR _25357_/D sky130_fd_sc_hd__and3_4
XFILLER_18_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14714_ _21403_/A VGND VGND VPWR VPWR _14714_/X sky130_fd_sc_hd__buf_2
X_17502_ _17605_/A VGND VGND VPWR VPWR _17600_/C sky130_fd_sc_hd__inv_2
X_11926_ _11947_/A VGND VGND VPWR VPWR _11926_/X sky130_fd_sc_hd__buf_2
X_18482_ _18482_/A _18482_/B VGND VGND VPWR VPWR _18483_/B sky130_fd_sc_hd__nor2_4
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20899__B2 _20886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15694_ _15693_/Y VGND VGND VPWR VPWR _15694_/X sky130_fd_sc_hd__buf_2
XANTENNA__24987__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17433_ _17431_/Y _17432_/X _16852_/X _17432_/X VGND VGND VPWR VPWR _17433_/X sky130_fd_sc_hd__a2bb2o_4
X_14645_ _14645_/A VGND VGND VPWR VPWR _18087_/A sky130_fd_sc_hd__inv_2
X_11857_ _11856_/X VGND VGND VPWR VPWR _15986_/A sky130_fd_sc_hd__buf_2
XANTENNA__24916__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17364_ _17363_/X VGND VGND VPWR VPWR _24336_/D sky130_fd_sc_hd__inv_2
X_14576_ _14554_/Y _14557_/X _14574_/X _25085_/Q _14575_/Y VGND VGND VPWR VPWR _25085_/D
+ sky130_fd_sc_hd__a32o_4
X_11788_ HWDATA[18] VGND VGND VPWR VPWR _11788_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_34_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_69_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16315_ _22899_/A VGND VGND VPWR VPWR _16315_/Y sky130_fd_sc_hd__inv_2
X_19103_ _19102_/Y _19098_/X _18919_/X _19098_/A VGND VGND VPWR VPWR _19103_/X sky130_fd_sc_hd__a2bb2o_4
X_13527_ _13514_/Y _13527_/B VGND VGND VPWR VPWR _13527_/X sky130_fd_sc_hd__and2_4
XANTENNA__15527__B1 HADDR[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_97_0_HCLK clkbuf_6_48_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_97_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17295_ _17295_/A _17295_/B VGND VGND VPWR VPWR _17295_/X sky130_fd_sc_hd__or2_4
X_19034_ _23869_/Q VGND VGND VPWR VPWR _19034_/Y sky130_fd_sc_hd__inv_2
X_16246_ _24643_/Q VGND VGND VPWR VPWR _16246_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13458_ _13426_/A _13458_/B VGND VGND VPWR VPWR _13458_/X sky130_fd_sc_hd__or2_4
XANTENNA__16036__A1_N _16033_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20928__A1_N _20909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12409_ _12389_/A _12409_/B _12408_/X VGND VGND VPWR VPWR _25447_/D sky130_fd_sc_hd__and3_4
X_16177_ _13739_/B _16176_/Y _14770_/B _16176_/Y VGND VGND VPWR VPWR _16177_/X sky130_fd_sc_hd__a2bb2o_4
X_13389_ _13421_/A _13387_/X _13389_/C VGND VGND VPWR VPWR _13389_/X sky130_fd_sc_hd__and3_4
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15128_ _24975_/Q VGND VGND VPWR VPWR _15128_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_3_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_126_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15674__A _16373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15059_ _15246_/A VGND VGND VPWR VPWR _15198_/A sky130_fd_sc_hd__buf_2
X_19936_ _19943_/A VGND VGND VPWR VPWR _19936_/X sky130_fd_sc_hd__buf_2
XFILLER_99_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18050__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19867_ _19866_/X VGND VGND VPWR VPWR _19880_/A sky130_fd_sc_hd__inv_2
XANTENNA__11707__A _24936_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18818_ _18799_/A _18818_/B _18817_/Y VGND VGND VPWR VPWR _24115_/D sky130_fd_sc_hd__and3_4
XFILLER_110_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19798_ _21375_/B _19793_/X _19797_/X _19793_/X VGND VGND VPWR VPWR _19798_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18749_ _18749_/A _18747_/A VGND VGND VPWR VPWR _18749_/X sky130_fd_sc_hd__or2_4
XFILLER_97_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21760_ _21247_/A VGND VGND VPWR VPWR _21763_/A sky130_fd_sc_hd__buf_2
X_20711_ _20711_/A VGND VGND VPWR VPWR _24004_/D sky130_fd_sc_hd__inv_2
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24657__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21691_ _21691_/A _22998_/A VGND VGND VPWR VPWR _21691_/X sky130_fd_sc_hd__or2_4
XANTENNA__16619__A1_N _16618_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23430_ _23478_/CLK _23430_/D VGND VGND VPWR VPWR _20268_/A sky130_fd_sc_hd__dfxtp_4
X_20642_ _20642_/A _20642_/B VGND VGND VPWR VPWR _20643_/B sky130_fd_sc_hd__nand2_4
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17507__A1 _25526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20573_ _20572_/X VGND VGND VPWR VPWR _23939_/D sky130_fd_sc_hd__inv_2
XANTENNA__15518__B1 HADDR[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23361_ _21004_/X VGND VGND VPWR VPWR IRQ[7] sky130_fd_sc_hd__buf_2
XFILLER_137_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25100_ _24077_/CLK _14499_/X HRESETn VGND VGND VPWR VPWR _23919_/D sky130_fd_sc_hd__dfrtp_4
X_22312_ _11990_/Y _12096_/X _11989_/Y _12071_/A VGND VGND VPWR VPWR _22312_/X sky130_fd_sc_hd__o22a_4
XFILLER_34_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23292_ _24564_/Q _23166_/X _23130_/X VGND VGND VPWR VPWR _23292_/X sky130_fd_sc_hd__o21a_4
X_25031_ _23989_/CLK _14867_/X HRESETn VGND VGND VPWR VPWR _25031_/Q sky130_fd_sc_hd__dfrtp_4
X_22243_ _22246_/A _22243_/B VGND VGND VPWR VPWR _22243_/X sky130_fd_sc_hd__or2_4
XANTENNA__22803__A2 _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22174_ _22174_/A VGND VGND VPWR VPWR _22174_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21586__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20490__A _20490_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25445__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21125_ _21119_/Y _21125_/B _21123_/X _21124_/X VGND VGND VPWR VPWR _21125_/X sky130_fd_sc_hd__and4_4
XANTENNA__19056__A _19055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22567__A1 _12944_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21056_ _21729_/A _21055_/Y _24700_/Q _21729_/A VGND VGND VPWR VPWR _21056_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18895__A _18895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23009__C _22812_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20007_ _20014_/A VGND VGND VPWR VPWR _20007_/X sky130_fd_sc_hd__buf_2
XFILLER_115_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24815_ _25330_/CLK _24815_/D HRESETn VGND VGND VPWR VPWR _24815_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12760_ _25376_/Q _12758_/Y _12747_/A _12759_/Y VGND VGND VPWR VPWR _12760_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24746_ _24766_/CLK _15974_/X HRESETn VGND VGND VPWR VPWR _24746_/Q sky130_fd_sc_hd__dfrtp_4
X_21958_ _21958_/A _19604_/Y VGND VGND VPWR VPWR _21958_/X sky130_fd_sc_hd__and2_4
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18943__B1 _17443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _12049_/A VGND VGND VPWR VPWR _15991_/A sky130_fd_sc_hd__buf_2
XFILLER_37_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _20909_/A VGND VGND VPWR VPWR _20909_/X sky130_fd_sc_hd__buf_2
XANTENNA__15757__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24398__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12691_/A VGND VGND VPWR VPWR _12691_/Y sky130_fd_sc_hd__inv_2
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24677_ _24673_/CLK _16145_/X HRESETn VGND VGND VPWR VPWR _22484_/A sky130_fd_sc_hd__dfrtp_4
X_21889_ _21885_/X _21889_/B _21888_/X VGND VGND VPWR VPWR _21889_/X sky130_fd_sc_hd__and3_4
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _25125_/Q VGND VGND VPWR VPWR _14430_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23628_ _23635_/CLK _23628_/D VGND VGND VPWR VPWR _23628_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15772__A3 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _14355_/X _14359_/X _12076_/A _14360_/X VGND VGND VPWR VPWR _25147_/D sky130_fd_sc_hd__o22a_4
XFILLER_35_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15509__B1 HADDR[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23559_ _25055_/CLK _19924_/X VGND VGND VPWR VPWR _19922_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16100_ _24694_/Q VGND VGND VPWR VPWR _16100_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _13312_/A _13312_/B VGND VGND VPWR VPWR _13313_/C sky130_fd_sc_hd__or2_4
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17080_ _17029_/A _17079_/X _17056_/X VGND VGND VPWR VPWR _17080_/Y sky130_fd_sc_hd__a21oi_4
X_14292_ _14292_/A VGND VGND VPWR VPWR _14292_/Y sky130_fd_sc_hd__inv_2
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16031_ _24720_/Q VGND VGND VPWR VPWR _16031_/Y sky130_fd_sc_hd__inv_2
X_13243_ _13188_/A _13240_/X _13243_/C VGND VGND VPWR VPWR _13243_/X sky130_fd_sc_hd__and3_4
X_25229_ _23967_/CLK _25229_/D HRESETn VGND VGND VPWR VPWR _14042_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_136_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12743__B1 _12842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13174_ _13173_/X VGND VGND VPWR VPWR _13174_/X sky130_fd_sc_hd__buf_2
XFILLER_124_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23962__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12125_ _12125_/A _24096_/Q VGND VGND VPWR VPWR _12126_/B sky130_fd_sc_hd__and2_4
XANTENNA__15494__A _15490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17982_ _17996_/A VGND VGND VPWR VPWR _17982_/X sky130_fd_sc_hd__buf_2
XFILLER_97_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22558__B2 _22922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25115__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19721_ _11856_/X VGND VGND VPWR VPWR _19721_/X sky130_fd_sc_hd__buf_2
X_12056_ _11725_/B VGND VGND VPWR VPWR _15652_/D sky130_fd_sc_hd__buf_2
X_16933_ _16133_/Y _17752_/A _16133_/Y _17752_/A VGND VGND VPWR VPWR _16933_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18226__A2 _18210_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15644__D _14433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19652_ _23655_/Q VGND VGND VPWR VPWR _19652_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16864_ _16862_/Y _16859_/X _16863_/X _16859_/X VGND VGND VPWR VPWR _24399_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18603_ _18603_/A VGND VGND VPWR VPWR _18603_/X sky130_fd_sc_hd__buf_2
X_15815_ _12341_/Y _15812_/X _11791_/X _15812_/X VGND VGND VPWR VPWR _24824_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22758__C _22736_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16795_ _16795_/A _16728_/B VGND VGND VPWR VPWR _16801_/A sky130_fd_sc_hd__nor2_4
X_19583_ _19582_/X VGND VGND VPWR VPWR _21364_/C sky130_fd_sc_hd__inv_2
XFILLER_92_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22120__A _21306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15746_ _15728_/X _15742_/X _15745_/X _24856_/Q _15740_/X VGND VGND VPWR VPWR _15746_/X
+ sky130_fd_sc_hd__a32o_4
X_18534_ _18405_/Y _18539_/B _18487_/X VGND VGND VPWR VPWR _18534_/Y sky130_fd_sc_hd__a21oi_4
X_12958_ _12957_/X VGND VGND VPWR VPWR _25363_/D sky130_fd_sc_hd__inv_2
XANTENNA__22730__A1 _17252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11909_ _11908_/X VGND VGND VPWR VPWR _11909_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24750__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15677_ _15677_/A VGND VGND VPWR VPWR _15677_/X sky130_fd_sc_hd__buf_2
X_18465_ _18420_/Y _18540_/A _18465_/C VGND VGND VPWR VPWR _18523_/A sky130_fd_sc_hd__or3_4
XFILLER_34_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15748__B1 _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12889_ _12889_/A VGND VGND VPWR VPWR _12890_/B sky130_fd_sc_hd__inv_2
XANTENNA__22774__B _22644_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14628_ _14628_/A VGND VGND VPWR VPWR _14628_/Y sky130_fd_sc_hd__inv_2
X_17416_ _17416_/A _14223_/B VGND VGND VPWR VPWR _17432_/A sky130_fd_sc_hd__nor2_4
XFILLER_53_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24068__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18396_ _18391_/X _18392_/X _18394_/X _18395_/X VGND VGND VPWR VPWR _18396_/X sky130_fd_sc_hd__or4_4
XANTENNA__14420__B1 _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17347_ _17245_/X _17347_/B VGND VGND VPWR VPWR _17348_/B sky130_fd_sc_hd__or2_4
XANTENNA__15669__A _15668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14559_ _14559_/A VGND VGND VPWR VPWR _14559_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22494__B1 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18045__A _18221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17278_ _17266_/A _17278_/B _17278_/C VGND VGND VPWR VPWR _17278_/X sky130_fd_sc_hd__and3_4
XANTENNA__22790__A _22790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_121_0_HCLK clkbuf_7_60_0_HCLK/X VGND VGND VPWR VPWR _24517_/CLK sky130_fd_sc_hd__clkbuf_1
X_16229_ _16227_/Y _16225_/X _16228_/X _16225_/X VGND VGND VPWR VPWR _16229_/X sky130_fd_sc_hd__a2bb2o_4
X_19017_ HWDATA[7] VGND VGND VPWR VPWR _19017_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_184_0_HCLK clkbuf_7_92_0_HCLK/X VGND VGND VPWR VPWR _23396_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22261__A3 _22256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21837__C _22695_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19919_ _19918_/Y _19916_/X _19787_/X _19916_/X VGND VGND VPWR VPWR _19919_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22949__B _22832_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22930_ _24452_/Q _22421_/X _22885_/X VGND VGND VPWR VPWR _22930_/X sky130_fd_sc_hd__o21a_4
XFILLER_25_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23126__A _23126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15987__B1 _15986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15851__B _15851_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24838__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22861_ _22770_/X _22860_/X _22479_/X _16029_/A _22480_/X VGND VGND VPWR VPWR _22861_/X
+ sky130_fd_sc_hd__a32o_4
X_24600_ _24600_/CLK _16364_/X HRESETn VGND VGND VPWR VPWR _24600_/Q sky130_fd_sc_hd__dfrtp_4
X_21812_ _21452_/A _21812_/B _21811_/X VGND VGND VPWR VPWR _21812_/X sky130_fd_sc_hd__and3_4
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22792_ _22792_/A _22791_/X VGND VGND VPWR VPWR _22792_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__17180__A2_N _17242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24531_ _24561_/CLK _16552_/X HRESETn VGND VGND VPWR VPWR _24531_/Q sky130_fd_sc_hd__dfrtp_4
X_21743_ _21103_/X _21741_/Y _21587_/X _21742_/X VGND VGND VPWR VPWR _21744_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24491__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24420__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24462_ _24462_/CLK _16735_/X HRESETn VGND VGND VPWR VPWR _15005_/A sky130_fd_sc_hd__dfrtp_4
X_21674_ _21484_/A _19527_/Y VGND VGND VPWR VPWR _21674_/X sky130_fd_sc_hd__or2_4
XFILLER_36_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23413_ _23533_/CLK _20314_/X VGND VGND VPWR VPWR _23413_/Q sky130_fd_sc_hd__dfxtp_4
X_20625_ _20625_/A _20624_/Y _20611_/C VGND VGND VPWR VPWR _20625_/X sky130_fd_sc_hd__and3_4
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14962__B2 _24416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24393_ _23846_/CLK _16889_/X HRESETn VGND VGND VPWR VPWR _19841_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19350__B1 _19349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23344_ _23344_/A _23344_/B VGND VGND VPWR VPWR _23344_/X sky130_fd_sc_hd__and2_4
X_20556_ _20556_/A VGND VGND VPWR VPWR _20556_/X sky130_fd_sc_hd__buf_2
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16164__B1 _15840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_80_0_HCLK clkbuf_7_81_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_80_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23275_ _24629_/Q _21519_/B VGND VGND VPWR VPWR _23275_/X sky130_fd_sc_hd__or2_4
X_20487_ _20487_/A _20486_/X VGND VGND VPWR VPWR _20487_/X sky130_fd_sc_hd__or2_4
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25014_ _25016_/CLK _25014_/D HRESETn VGND VGND VPWR VPWR _25014_/Q sky130_fd_sc_hd__dfrtp_4
X_22226_ _22229_/A _22226_/B VGND VGND VPWR VPWR _22226_/X sky130_fd_sc_hd__or2_4
XFILLER_133_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22157_ _16451_/A _22154_/X _22157_/C VGND VGND VPWR VPWR _22157_/X sky130_fd_sc_hd__and3_4
XFILLER_105_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21108_ _15638_/Y _21108_/B VGND VGND VPWR VPWR _21108_/X sky130_fd_sc_hd__or2_4
XFILLER_43_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22088_ _22088_/A VGND VGND VPWR VPWR _22701_/A sky130_fd_sc_hd__buf_2
XFILLER_94_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13930_ _13930_/A _13930_/B _13942_/C _13930_/D VGND VGND VPWR VPWR _13931_/A sky130_fd_sc_hd__or4_4
XFILLER_75_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21039_ _21029_/X _21035_/X _22664_/B _21038_/X VGND VGND VPWR VPWR _21040_/C sky130_fd_sc_hd__a211o_4
XFILLER_86_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13861_ _13860_/X VGND VGND VPWR VPWR _13861_/X sky130_fd_sc_hd__buf_2
XANTENNA__24579__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15600_ _15588_/A VGND VGND VPWR VPWR _15600_/X sky130_fd_sc_hd__buf_2
X_12812_ _12926_/A VGND VGND VPWR VPWR _12849_/A sky130_fd_sc_hd__inv_2
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16580_ _16579_/Y _16575_/X _16410_/X _16575_/X VGND VGND VPWR VPWR _16580_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24508__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13792_ _13791_/X VGND VGND VPWR VPWR _21996_/A sky130_fd_sc_hd__inv_2
XANTENNA__14377__B _14377_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15531_ _11726_/B VGND VGND VPWR VPWR _15531_/Y sky130_fd_sc_hd__inv_2
X_12743_ _12842_/A _24783_/Q _12842_/A _24783_/Q VGND VGND VPWR VPWR _12743_/X sky130_fd_sc_hd__a2bb2o_4
X_24729_ _24345_/CLK _24729_/D HRESETn VGND VGND VPWR VPWR _24729_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17195__A2 _23246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18250_ _11661_/Y _18249_/X _17421_/X _18249_/X VGND VGND VPWR VPWR _24219_/D sky130_fd_sc_hd__a2bb2o_4
X_15462_ _15462_/A _14223_/B VGND VGND VPWR VPWR _15476_/A sky130_fd_sc_hd__nor2_4
XANTENNA__24161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12674_ _12567_/Y _12674_/B VGND VGND VPWR VPWR _12674_/X sky130_fd_sc_hd__or2_4
XFILLER_54_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17193_/X _17201_/B _17201_/C _17201_/D VGND VGND VPWR VPWR _17202_/D sky130_fd_sc_hd__or4_4
XFILLER_93_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ HWDATA[6] VGND VGND VPWR VPWR _15623_/A sky130_fd_sc_hd__buf_2
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18181_ _18181_/A _18181_/B _18181_/C VGND VGND VPWR VPWR _18185_/B sky130_fd_sc_hd__and3_4
XANTENNA__15489__A _24064_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _15299_/B _15392_/X VGND VGND VPWR VPWR _15400_/B sky130_fd_sc_hd__or2_4
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17132_ _17038_/C _17148_/A VGND VGND VPWR VPWR _17132_/X sky130_fd_sc_hd__or2_4
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14344_ _14348_/A VGND VGND VPWR VPWR _14344_/X sky130_fd_sc_hd__buf_2
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16155__B1 _16064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17063_ _16981_/Y _17061_/A VGND VGND VPWR VPWR _17063_/X sky130_fd_sc_hd__or2_4
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25367__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14275_ _25172_/Q VGND VGND VPWR VPWR _14275_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15902__B1 _15620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16014_ _24727_/Q VGND VGND VPWR VPWR _16014_/Y sky130_fd_sc_hd__inv_2
X_13226_ _13310_/A _18927_/A VGND VGND VPWR VPWR _13226_/X sky130_fd_sc_hd__or2_4
XANTENNA__22779__B2 _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12192__B2 _24761_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13157_ _13156_/X VGND VGND VPWR VPWR _13188_/A sky130_fd_sc_hd__buf_2
XANTENNA__16113__A _16094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12108_ _12106_/Y _12102_/X _11833_/X _12107_/X VGND VGND VPWR VPWR _25463_/D sky130_fd_sc_hd__a2bb2o_4
X_13088_ _12292_/Y _13087_/X _13031_/X VGND VGND VPWR VPWR _13088_/Y sky130_fd_sc_hd__a21oi_4
X_17965_ _14645_/A VGND VGND VPWR VPWR _18176_/A sky130_fd_sc_hd__buf_2
XFILLER_100_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19704_ _23636_/Q VGND VGND VPWR VPWR _19704_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15952__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12039_ _12038_/Y _12034_/X _12040_/A _12034_/X VGND VGND VPWR VPWR _25478_/D sky130_fd_sc_hd__a2bb2o_4
X_16916_ _16916_/A VGND VGND VPWR VPWR _16916_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19424__A _19423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21535__A1_N _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17896_ _17893_/Y _17889_/X _17895_/Y VGND VGND VPWR VPWR _17896_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19635_ _21177_/B _19628_/X _19488_/X _19628_/A VGND VGND VPWR VPWR _23661_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16847_ _24405_/Q VGND VGND VPWR VPWR _16847_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24931__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13472__A _11867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24249__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19566_ _23682_/Q VGND VGND VPWR VPWR _22023_/B sky130_fd_sc_hd__inv_2
XFILLER_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16778_ _16773_/A VGND VGND VPWR VPWR _16778_/X sky130_fd_sc_hd__buf_2
XFILLER_59_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_5_23_0_HCLK_A clkbuf_5_22_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15984__A3 _15836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18517_ _18517_/A _18517_/B _18516_/X VGND VGND VPWR VPWR _18517_/X sky130_fd_sc_hd__and3_4
X_15729_ HWDATA[23] VGND VGND VPWR VPWR _15729_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19497_ _23707_/Q VGND VGND VPWR VPWR _22249_/B sky130_fd_sc_hd__inv_2
XANTENNA__16783__A _16733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18448_ _16253_/Y _18393_/A _16261_/Y _24148_/Q VGND VGND VPWR VPWR _18448_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17591__C1 _17590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18379_ _24182_/Q VGND VGND VPWR VPWR _18379_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11720__A _16371_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20410_ _20409_/Y _20405_/X _15768_/X _20405_/X VGND VGND VPWR VPWR _23374_/D sky130_fd_sc_hd__a2bb2o_4
X_21390_ _21393_/A _19925_/Y VGND VGND VPWR VPWR _21390_/X sky130_fd_sc_hd__or2_4
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16925__A2_N _17758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20341_ _22332_/B _20340_/X _19612_/A _20340_/X VGND VGND VPWR VPWR _20341_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18503__A _18503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25037__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20272_ _20996_/B _14796_/C VGND VGND VPWR VPWR _20272_/X sky130_fd_sc_hd__or2_4
X_23060_ _24525_/Q _22922_/X _22923_/X _23059_/X VGND VGND VPWR VPWR _23061_/C sky130_fd_sc_hd__a211o_4
XANTENNA__14750__B _14744_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22011_ _21671_/A _22011_/B _22010_/X VGND VGND VPWR VPWR _22011_/X sky130_fd_sc_hd__and3_4
XANTENNA__21442__A1 _12976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21864__A _22664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15862__A _15702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23962_ _24070_/CLK _20999_/X HRESETn VGND VGND VPWR VPWR _23962_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22913_ _22913_/A VGND VGND VPWR VPWR _22914_/B sky130_fd_sc_hd__buf_2
XANTENNA__24672__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23893_ _23905_/CLK _23893_/D VGND VGND VPWR VPWR _18965_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_83_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15424__A2 _15316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16621__B2 _16545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24601__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22844_ _23034_/A VGND VGND VPWR VPWR _22844_/X sky130_fd_sc_hd__buf_2
XANTENNA__22695__A _24447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22775_ _15544_/X VGND VGND VPWR VPWR _22775_/X sky130_fd_sc_hd__buf_2
XFILLER_25_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24514_ _24517_/CLK _16593_/X HRESETn VGND VGND VPWR VPWR _16592_/A sky130_fd_sc_hd__dfrtp_4
X_21726_ _21560_/X _21724_/X _21566_/X _21725_/X VGND VGND VPWR VPWR _21727_/A sky130_fd_sc_hd__o22a_4
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16385__B1 _16384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25494_ _23714_/CLK _25494_/D HRESETn VGND VGND VPWR VPWR _11937_/A sky130_fd_sc_hd__dfrtp_4
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21104__A _15551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24445_ _24462_/CLK _16768_/X HRESETn VGND VGND VPWR VPWR _24445_/Q sky130_fd_sc_hd__dfrtp_4
X_21657_ _21465_/A _19963_/Y VGND VGND VPWR VPWR _21659_/B sky130_fd_sc_hd__or2_4
XFILLER_32_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19323__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20608_ _20607_/X VGND VGND VPWR VPWR _20608_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12390_ _12382_/X _12390_/B VGND VGND VPWR VPWR _12391_/B sky130_fd_sc_hd__and2_4
XFILLER_21_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24376_ _24376_/CLK _17112_/X HRESETn VGND VGND VPWR VPWR _17030_/A sky130_fd_sc_hd__dfrtp_4
X_21588_ _21581_/X VGND VGND VPWR VPWR _21588_/X sky130_fd_sc_hd__buf_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25460__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23327_ _24598_/Q _23327_/B VGND VGND VPWR VPWR _23327_/X sky130_fd_sc_hd__or2_4
X_20539_ _20539_/A _20537_/Y _20558_/C VGND VGND VPWR VPWR _20539_/X sky130_fd_sc_hd__and3_4
X_14060_ _14052_/X _14076_/A VGND VGND VPWR VPWR _14060_/X sky130_fd_sc_hd__or2_4
XFILLER_84_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23258_ _14930_/A _21533_/X _22090_/X _23257_/X VGND VGND VPWR VPWR _23259_/C sky130_fd_sc_hd__a211o_4
XFILLER_4_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13011_ _13011_/A VGND VGND VPWR VPWR _13011_/Y sky130_fd_sc_hd__inv_2
X_22209_ _22193_/X _22209_/B VGND VGND VPWR VPWR _22209_/X sky130_fd_sc_hd__or2_4
XANTENNA__17637__B1 _17590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13557__A _13557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23189_ _23105_/X _23186_/Y _23150_/X _23188_/X VGND VGND VPWR VPWR _23189_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_24_0_HCLK clkbuf_7_12_0_HCLK/X VGND VGND VPWR VPWR _25478_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_87_0_HCLK clkbuf_8_87_0_HCLK/A VGND VGND VPWR VPWR _24950_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16868__A _16880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14962_ _14961_/X _24416_/Q _14960_/Y _24416_/Q VGND VGND VPWR VPWR _14962_/X sky130_fd_sc_hd__a2bb2o_4
X_17750_ _16918_/Y _17846_/A _16898_/A _17750_/D VGND VGND VPWR VPWR _17750_/X sky130_fd_sc_hd__or4_4
XFILLER_82_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16701_ _16699_/Y _16695_/X _16604_/X _16700_/X VGND VGND VPWR VPWR _24474_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13913_ _13927_/A VGND VGND VPWR VPWR _13913_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14893_ _25020_/Q VGND VGND VPWR VPWR _14893_/Y sky130_fd_sc_hd__inv_2
X_17681_ _17624_/A VGND VGND VPWR VPWR _17681_/X sky130_fd_sc_hd__buf_2
X_19420_ _17442_/X VGND VGND VPWR VPWR _19420_/X sky130_fd_sc_hd__buf_2
X_13844_ _13572_/Y _13839_/X _13800_/X _13843_/X VGND VGND VPWR VPWR _25245_/D sky130_fd_sc_hd__a2bb2o_4
X_16632_ _16631_/X VGND VGND VPWR VPWR _16632_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24342__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19351_ _18214_/B VGND VGND VPWR VPWR _19351_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13775_ _13774_/Y VGND VGND VPWR VPWR _13775_/X sky130_fd_sc_hd__buf_2
X_16563_ _16558_/A VGND VGND VPWR VPWR _16563_/X sky130_fd_sc_hd__buf_2
X_18302_ _18299_/X _18301_/X _18296_/X VGND VGND VPWR VPWR _18302_/X sky130_fd_sc_hd__o21a_4
X_12726_ _12616_/B _12702_/X _12724_/B _12653_/X VGND VGND VPWR VPWR _12726_/X sky130_fd_sc_hd__a211o_4
X_15514_ _15513_/Y _15511_/X HADDR[13] _15511_/X VGND VGND VPWR VPWR _15514_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16494_ _16493_/Y _16491_/X _16408_/X _16491_/X VGND VGND VPWR VPWR _16494_/X sky130_fd_sc_hd__a2bb2o_4
X_19282_ _23781_/Q VGND VGND VPWR VPWR _21235_/B sky130_fd_sc_hd__inv_2
XFILLER_95_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15445_ _13920_/X _15437_/X _15432_/X _13919_/X _15444_/X VGND VGND VPWR VPWR _15445_/X
+ sky130_fd_sc_hd__a32o_4
X_18233_ _18233_/A VGND VGND VPWR VPWR _18233_/X sky130_fd_sc_hd__buf_2
XFILLER_19_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12657_ _12657_/A _12652_/X _12656_/Y VGND VGND VPWR VPWR _12657_/X sky130_fd_sc_hd__and3_4
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19314__B1 _19313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15376_ _15130_/Y _15352_/B _15318_/A _15373_/Y VGND VGND VPWR VPWR _15376_/X sky130_fd_sc_hd__a211o_4
X_18164_ _18196_/A _18164_/B VGND VGND VPWR VPWR _18164_/X sky130_fd_sc_hd__or2_4
X_12588_ _25410_/Q _12586_/Y _12611_/B _24862_/Q VGND VGND VPWR VPWR _12588_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14327_ _14327_/A VGND VGND VPWR VPWR _14327_/Y sky130_fd_sc_hd__inv_2
X_17115_ _17108_/A _17105_/B _17115_/C VGND VGND VPWR VPWR _24375_/D sky130_fd_sc_hd__and3_4
X_18095_ _18191_/A _18095_/B _18094_/X VGND VGND VPWR VPWR _18095_/X sky130_fd_sc_hd__and3_4
X_17046_ _17036_/Y _17120_/A _17045_/X VGND VGND VPWR VPWR _17091_/B sky130_fd_sc_hd__or3_4
X_14258_ _14258_/A _14223_/B VGND VGND VPWR VPWR _14271_/A sky130_fd_sc_hd__nor2_4
XFILLER_131_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13209_ _24190_/Q VGND VGND VPWR VPWR _13225_/A sky130_fd_sc_hd__buf_2
X_14189_ _15991_/A _11719_/B _15991_/C _16369_/D VGND VGND VPWR VPWR _14190_/B sky130_fd_sc_hd__or4_4
XFILLER_112_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18997_ _18996_/X VGND VGND VPWR VPWR _18997_/X sky130_fd_sc_hd__buf_2
XFILLER_61_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17948_ _17955_/A _19309_/A VGND VGND VPWR VPWR _17950_/B sky130_fd_sc_hd__or2_4
XFILLER_39_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17879_ _17748_/Y _17878_/X _16955_/X VGND VGND VPWR VPWR _17879_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_96_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18993__A _19642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19618_ _19618_/A VGND VGND VPWR VPWR _19618_/X sky130_fd_sc_hd__buf_2
XANTENNA__11715__A _11714_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20890_ _20888_/Y _20884_/Y _20889_/X VGND VGND VPWR VPWR _20890_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24012__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19549_ _23688_/Q VGND VGND VPWR VPWR _19549_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22152__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22560_ _22560_/A _22598_/B VGND VGND VPWR VPWR _22560_/X sky130_fd_sc_hd__and2_4
XFILLER_62_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16367__B1 _16366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21511_ _21069_/A VGND VGND VPWR VPWR _21511_/X sky130_fd_sc_hd__buf_2
X_22491_ _17350_/A _22424_/A _12954_/A _22288_/X VGND VGND VPWR VPWR _22492_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19305__B1 _19191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24230_ _23826_/CLK _24230_/D HRESETn VGND VGND VPWR VPWR _24230_/Q sky130_fd_sc_hd__dfrtp_4
X_21442_ _12976_/A _21438_/X _21441_/X VGND VGND VPWR VPWR _21442_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16119__B1 _15959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24161_ _24162_/CLK _24161_/D HRESETn VGND VGND VPWR VPWR _18461_/A sky130_fd_sc_hd__dfrtp_4
X_21373_ _21393_/A _21373_/B VGND VGND VPWR VPWR _21374_/C sky130_fd_sc_hd__or2_4
XFILLER_68_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23112_ _22975_/X _23110_/X _23044_/X _11763_/A _23111_/X VGND VGND VPWR VPWR _23112_/X
+ sky130_fd_sc_hd__a32o_4
X_20324_ _20317_/X _19586_/D _11842_/A _21978_/C _20326_/A VGND VGND VPWR VPWR _20324_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24092_ _25246_/CLK _12026_/C HRESETn VGND VGND VPWR VPWR _12020_/A sky130_fd_sc_hd__dfrtp_4
X_23043_ _23043_/A _22864_/X VGND VGND VPWR VPWR _23043_/X sky130_fd_sc_hd__or2_4
X_20255_ _22367_/B _20254_/X _19777_/A _20254_/X VGND VGND VPWR VPWR _23436_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_240_0_HCLK clkbuf_8_241_0_HCLK/A VGND VGND VPWR VPWR _24018_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20186_ _20186_/A VGND VGND VPWR VPWR _20186_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24853__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16688__A _16664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24994_ _24984_/CLK _15314_/X HRESETn VGND VGND VPWR VPWR _24994_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23945_ _25199_/CLK scl_i_S4 HRESETn VGND VGND VPWR VPWR _23945_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11890_ _11874_/Y _11887_/X _25506_/Q _11889_/Y VGND VGND VPWR VPWR _25506_/D sky130_fd_sc_hd__o22a_4
X_23876_ _25485_/CLK _19019_/X VGND VGND VPWR VPWR _23876_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15948__A3 HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22827_ _22827_/A VGND VGND VPWR VPWR _22827_/X sky130_fd_sc_hd__buf_2
XANTENNA__13840__A _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13560_ _25081_/Q VGND VGND VPWR VPWR _14572_/A sky130_fd_sc_hd__inv_2
XFILLER_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22758_ _22725_/X _22732_/Y _22736_/X _22758_/D VGND VGND VPWR VPWR HRDATA[15] sky130_fd_sc_hd__or4_4
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12511_ _12510_/Y _24853_/Q _12510_/Y _24853_/Q VGND VGND VPWR VPWR _12511_/X sky130_fd_sc_hd__a2bb2o_4
X_21709_ _21709_/A _22111_/B VGND VGND VPWR VPWR _21709_/Y sky130_fd_sc_hd__nand2_4
X_13491_ _25305_/Q VGND VGND VPWR VPWR _13491_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25477_ _25461_/CLK _25477_/D HRESETn VGND VGND VPWR VPWR _12040_/A sky130_fd_sc_hd__dfrtp_4
X_22689_ _24227_/Q _22613_/B VGND VGND VPWR VPWR _22689_/Y sky130_fd_sc_hd__nor2_4
X_15230_ _15230_/A VGND VGND VPWR VPWR _15230_/Y sky130_fd_sc_hd__inv_2
X_12442_ _12286_/C _12440_/X _12441_/Y VGND VGND VPWR VPWR _25439_/D sky130_fd_sc_hd__o21a_4
XFILLER_60_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24428_ _24431_/CLK _16805_/X HRESETn VGND VGND VPWR VPWR _14905_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12395__A1 _12266_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15161_ _15154_/X _15161_/B _15161_/C _15160_/X VGND VGND VPWR VPWR _15161_/X sky130_fd_sc_hd__or4_4
X_12373_ _12378_/A _24810_/Q _25323_/Q _12344_/Y VGND VGND VPWR VPWR _12373_/X sky130_fd_sc_hd__a2bb2o_4
X_24359_ _24355_/CLK _17266_/X HRESETn VGND VGND VPWR VPWR _24359_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_50_0_HCLK clkbuf_6_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14112_ _25210_/Q VGND VGND VPWR VPWR _14119_/A sky130_fd_sc_hd__inv_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15092_ _24963_/Q VGND VGND VPWR VPWR _15092_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14043_ _14043_/A VGND VGND VPWR VPWR _14043_/Y sky130_fd_sc_hd__inv_2
X_18920_ _18918_/Y _18914_/X _18919_/X _18901_/Y VGND VGND VPWR VPWR _23909_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13287__A _13227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17982__A _17996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22603__B1 _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18851_ _16490_/Y _24132_/Q _16490_/Y _24132_/Q VGND VGND VPWR VPWR _18854_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24594__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20090__B1 _20089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17802_ _24268_/Q _17805_/B VGND VGND VPWR VPWR _17802_/X sky130_fd_sc_hd__or2_4
XFILLER_132_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24523__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18782_ _18782_/A VGND VGND VPWR VPWR _18782_/X sky130_fd_sc_hd__buf_2
X_15994_ _22915_/A _15993_/Y VGND VGND VPWR VPWR _15995_/A sky130_fd_sc_hd__and2_4
XFILLER_48_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17733_ _17733_/A _18318_/B _17726_/X _17733_/D VGND VGND VPWR VPWR _17734_/A sky130_fd_sc_hd__or4_4
X_14945_ _14945_/A VGND VGND VPWR VPWR _14945_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15652__D _15652_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17664_ _17528_/Y _17683_/A VGND VGND VPWR VPWR _17685_/A sky130_fd_sc_hd__or2_4
X_14876_ _14876_/A VGND VGND VPWR VPWR _14876_/Y sky130_fd_sc_hd__inv_2
X_19403_ _23739_/Q VGND VGND VPWR VPWR _19403_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16615_ _16613_/Y _16609_/X _16355_/X _16614_/X VGND VGND VPWR VPWR _16615_/X sky130_fd_sc_hd__a2bb2o_4
X_13827_ _22612_/A _13825_/X _11813_/X _13825_/X VGND VGND VPWR VPWR _13827_/X sky130_fd_sc_hd__a2bb2o_4
X_17595_ _17597_/B VGND VGND VPWR VPWR _17596_/B sky130_fd_sc_hd__inv_2
XANTENNA__18338__A1 _21504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19334_ _19333_/Y VGND VGND VPWR VPWR _19334_/X sky130_fd_sc_hd__buf_2
X_13758_ _13754_/A _13758_/B VGND VGND VPWR VPWR _13759_/A sky130_fd_sc_hd__and2_4
X_16546_ _16541_/Y _16545_/X _16376_/X _16545_/X VGND VGND VPWR VPWR _16546_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20145__B2 _20140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12709_ _12712_/A _12712_/B VGND VGND VPWR VPWR _12713_/B sky130_fd_sc_hd__or2_4
XANTENNA__25382__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19265_ _19264_/X VGND VGND VPWR VPWR _19278_/A sky130_fd_sc_hd__inv_2
XFILLER_56_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11830__B1 _11829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13689_ _13689_/A _13689_/B VGND VGND VPWR VPWR _13689_/X sky130_fd_sc_hd__or2_4
X_16477_ _16476_/Y _16474_/X _16300_/X _16474_/X VGND VGND VPWR VPWR _16477_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18216_ _18184_/A _18214_/X _18216_/C VGND VGND VPWR VPWR _18217_/C sky130_fd_sc_hd__and3_4
XANTENNA__25311__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15428_ _15428_/A _15427_/Y VGND VGND VPWR VPWR _15429_/B sky130_fd_sc_hd__or2_4
XFILLER_31_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19196_ _19014_/B _19038_/C _19038_/D _19038_/A VGND VGND VPWR VPWR _19197_/A sky130_fd_sc_hd__and4_4
XANTENNA__11701__C _11700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15359_ _15359_/A VGND VGND VPWR VPWR _15359_/Y sky130_fd_sc_hd__inv_2
X_18147_ _18080_/A _19029_/A VGND VGND VPWR VPWR _18149_/B sky130_fd_sc_hd__or2_4
XANTENNA__18053__A _18184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18078_ _17928_/X _18078_/B _18078_/C VGND VGND VPWR VPWR _18078_/X sky130_fd_sc_hd__and3_4
XFILLER_105_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17029_ _17029_/A _16976_/Y VGND VGND VPWR VPWR _17029_/X sky130_fd_sc_hd__or2_4
XFILLER_67_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20040_ _20040_/A VGND VGND VPWR VPWR _20040_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24264__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_70_0_HCLK clkbuf_8_71_0_HCLK/A VGND VGND VPWR VPWR _23978_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_100_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21991_ _17887_/Y _21977_/B VGND VGND VPWR VPWR _21991_/X sky130_fd_sc_hd__and2_4
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15536__A1_N _12059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23730_ _23718_/CLK _19432_/X VGND VGND VPWR VPWR _18034_/B sky130_fd_sc_hd__dfxtp_4
X_20942_ _20943_/A VGND VGND VPWR VPWR _20942_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _23396_/CLK _23661_/D VGND VGND VPWR VPWR _23661_/Q sky130_fd_sc_hd__dfxtp_4
X_20873_ _13663_/A VGND VGND VPWR VPWR _20873_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17547__A2_N _24308_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19526__B1 _11948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25400_ _25400_/CLK _12700_/Y HRESETn VGND VGND VPWR VPWR _12565_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17132__A _17038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22612_ _22612_/A _22726_/B VGND VGND VPWR VPWR _22612_/X sky130_fd_sc_hd__and2_4
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23592_ _23581_/CLK _19834_/X VGND VGND VPWR VPWR _19833_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25331_ _25351_/CLK _25331_/D HRESETn VGND VGND VPWR VPWR _12330_/A sky130_fd_sc_hd__dfrtp_4
X_22543_ _22736_/A _22539_/X _22543_/C VGND VGND VPWR VPWR _22543_/X sky130_fd_sc_hd__and3_4
XANTENNA__25052__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25262_ _25246_/CLK _13798_/X HRESETn VGND VGND VPWR VPWR _13786_/A sky130_fd_sc_hd__dfrtp_4
X_22474_ _22287_/A _22473_/X VGND VGND VPWR VPWR _22488_/C sky130_fd_sc_hd__and2_4
XANTENNA__16760__B1 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24213_ _24219_/CLK _24213_/D HRESETn VGND VGND VPWR VPWR _24213_/Q sky130_fd_sc_hd__dfrtp_4
X_21425_ _21525_/A VGND VGND VPWR VPWR _22998_/A sky130_fd_sc_hd__buf_2
X_25193_ _23989_/CLK _14208_/X HRESETn VGND VGND VPWR VPWR _14207_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_120_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24144_ _24133_/CLK _24144_/D HRESETn VGND VGND VPWR VPWR _24144_/Q sky130_fd_sc_hd__dfrtp_4
X_21356_ _21354_/Y _21143_/X _17434_/Y _21549_/B VGND VGND VPWR VPWR _21359_/C sky130_fd_sc_hd__o22a_4
XANTENNA__16512__B1 _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20307_ _21935_/B _20304_/X _19985_/X _20304_/X VGND VGND VPWR VPWR _23416_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24075_ _24117_/CLK _20494_/X HRESETn VGND VGND VPWR VPWR _24075_/Q sky130_fd_sc_hd__dfrtp_4
X_21287_ _22824_/A VGND VGND VPWR VPWR _21287_/Y sky130_fd_sc_hd__inv_2
X_23026_ _16110_/Y _22513_/B _22843_/X _11773_/Y _22846_/X VGND VGND VPWR VPWR _23026_/X
+ sky130_fd_sc_hd__o32a_4
X_20238_ _20232_/Y VGND VGND VPWR VPWR _20238_/X sky130_fd_sc_hd__buf_2
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13835__A _13835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17307__A _22659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20169_ _20169_/A VGND VGND VPWR VPWR _20182_/A sky130_fd_sc_hd__inv_2
XANTENNA__23010__B1 _21050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12991_ _13092_/A _12991_/B _13096_/A _12377_/Y VGND VGND VPWR VPWR _12991_/X sky130_fd_sc_hd__or4_4
XFILLER_131_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24977_ _24977_/CLK _24977_/D HRESETn VGND VGND VPWR VPWR _24977_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11942_ _11948_/A VGND VGND VPWR VPWR _11942_/Y sky130_fd_sc_hd__inv_2
X_14730_ _14727_/Y _14708_/X _14729_/Y VGND VGND VPWR VPWR _14730_/Y sky130_fd_sc_hd__o21ai_4
X_23928_ _25199_/CLK _20975_/X HRESETn VGND VGND VPWR VPWR _20976_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__20668__A _20664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14661_ _14661_/A VGND VGND VPWR VPWR _19038_/C sky130_fd_sc_hd__buf_2
XANTENNA__23044__A _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11873_ _11900_/A _11872_/X VGND VGND VPWR VPWR _11873_/X sky130_fd_sc_hd__or2_4
X_23859_ _23441_/CLK _23859_/D VGND VGND VPWR VPWR _13204_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18138__A _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13612_ _17929_/A VGND VGND VPWR VPWR _14641_/B sky130_fd_sc_hd__buf_2
X_16400_ _16389_/A VGND VGND VPWR VPWR _16400_/X sky130_fd_sc_hd__buf_2
XFILLER_72_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14592_ _14592_/A _14592_/B VGND VGND VPWR VPWR _14592_/Y sky130_fd_sc_hd__nand2_4
X_17380_ _17199_/Y _17377_/B VGND VGND VPWR VPWR _17380_/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22883__A _23170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13543_ _25247_/Q VGND VGND VPWR VPWR _13543_/Y sky130_fd_sc_hd__inv_2
X_16331_ _16329_/Y _16324_/X _16231_/X _16330_/X VGND VGND VPWR VPWR _24613_/D sky130_fd_sc_hd__a2bb2o_4
X_25529_ _24759_/CLK _11775_/X HRESETn VGND VGND VPWR VPWR _25529_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16262_ _16261_/Y _16259_/X _15474_/X _16259_/X VGND VGND VPWR VPWR _16262_/X sky130_fd_sc_hd__a2bb2o_4
X_19050_ _19049_/Y _19045_/X _18977_/X _19045_/X VGND VGND VPWR VPWR _23864_/D sky130_fd_sc_hd__a2bb2o_4
X_13474_ _25311_/Q VGND VGND VPWR VPWR _13474_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16751__B1 _16403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15213_ _15212_/X VGND VGND VPWR VPWR _15214_/B sky130_fd_sc_hd__inv_2
X_18001_ _18088_/A VGND VGND VPWR VPWR _18221_/A sky130_fd_sc_hd__buf_2
XFILLER_9_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12425_ _12389_/A _12415_/X _12425_/C VGND VGND VPWR VPWR _12425_/X sky130_fd_sc_hd__and3_4
XFILLER_12_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16193_ _16217_/A VGND VGND VPWR VPWR _16193_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15144_ _15144_/A VGND VGND VPWR VPWR _15389_/A sky130_fd_sc_hd__inv_2
X_12356_ _25339_/Q VGND VGND VPWR VPWR _13061_/A sky130_fd_sc_hd__inv_2
XANTENNA__24775__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15075_ _24994_/Q VGND VGND VPWR VPWR _15313_/A sky130_fd_sc_hd__inv_2
X_19952_ _19964_/A VGND VGND VPWR VPWR _19952_/X sky130_fd_sc_hd__buf_2
XFILLER_138_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12287_ _12242_/A _12235_/A _12285_/X _12432_/A VGND VGND VPWR VPWR _12287_/X sky130_fd_sc_hd__or4_4
XANTENNA__24704__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14026_ _14026_/A VGND VGND VPWR VPWR _14026_/Y sky130_fd_sc_hd__inv_2
X_18903_ _22363_/B _18902_/X _16863_/X _18902_/X VGND VGND VPWR VPWR _18903_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18256__B1 _16852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19883_ _19882_/Y _19880_/X _19632_/X _19880_/X VGND VGND VPWR VPWR _19883_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22123__A _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18834_ _24550_/Q _24129_/Q _16497_/Y _18753_/C VGND VGND VPWR VPWR _18838_/A sky130_fd_sc_hd__o22a_4
XFILLER_68_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13745__A _14705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12540__B2 _12539_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_57_0_HCLK clkbuf_6_28_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18765_ _18765_/A _18765_/B VGND VGND VPWR VPWR _18765_/X sky130_fd_sc_hd__or2_4
X_15977_ _12221_/Y _15975_/X _15756_/X _15975_/X VGND VGND VPWR VPWR _24744_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19756__B1 _19755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17716_ _21663_/A VGND VGND VPWR VPWR _17717_/A sky130_fd_sc_hd__buf_2
X_14928_ _25014_/Q _14927_/A _14926_/X _14927_/Y VGND VGND VPWR VPWR _14939_/A sky130_fd_sc_hd__o22a_4
X_18696_ _18696_/A _18695_/X VGND VGND VPWR VPWR _18704_/A sky130_fd_sc_hd__or2_4
XFILLER_58_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17647_ _17635_/B VGND VGND VPWR VPWR _17648_/B sky130_fd_sc_hd__inv_2
X_14859_ _14858_/X VGND VGND VPWR VPWR _14859_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17578_ _17528_/Y _17576_/Y _17578_/C _17577_/Y VGND VGND VPWR VPWR _17579_/C sky130_fd_sc_hd__or4_4
XFILLER_95_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19317_ _19317_/A VGND VGND VPWR VPWR _19317_/Y sky130_fd_sc_hd__inv_2
X_16529_ _16527_/Y _16524_/X _16528_/X _16524_/X VGND VGND VPWR VPWR _16529_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19248_ _23794_/Q VGND VGND VPWR VPWR _19248_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16742__B1 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12359__B2 _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19179_ _19178_/Y _19176_/X _19133_/X _19176_/X VGND VGND VPWR VPWR _19179_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21210_ _22824_/A VGND VGND VPWR VPWR _22790_/A sky130_fd_sc_hd__buf_2
XANTENNA__21094__A2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22291__A1 _25361_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22190_ _21240_/X _20047_/Y VGND VGND VPWR VPWR _22191_/C sky130_fd_sc_hd__or2_4
X_21141_ _21140_/Y _21335_/A _14881_/Y _14433_/A VGND VGND VPWR VPWR _21141_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24445__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21072_ _22464_/A VGND VGND VPWR VPWR _21073_/B sky130_fd_sc_hd__buf_2
XFILLER_120_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20023_ _20023_/A VGND VGND VPWR VPWR _20036_/A sky130_fd_sc_hd__inv_2
XFILLER_101_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17127__A _17023_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24900_ _24868_/CLK _15589_/X HRESETn VGND VGND VPWR VPWR _15587_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16031__A _24720_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22968__A _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21872__A _21009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15475__A1_N _15473_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24831_ _24852_/CLK _15806_/X HRESETn VGND VGND VPWR VPWR _24831_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15481__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12295__B1 _12294_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24762_ _25374_/CLK _15946_/X HRESETn VGND VGND VPWR VPWR _23178_/A sky130_fd_sc_hd__dfrtp_4
X_21974_ _18359_/Y _20329_/A _24188_/Q _20331_/Y VGND VGND VPWR VPWR _21974_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20357__B2 _20339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23713_ _24926_/CLK _23713_/D VGND VGND VPWR VPWR _23713_/Q sky130_fd_sc_hd__dfxtp_4
X_20925_ _24054_/Q VGND VGND VPWR VPWR _20925_/Y sky130_fd_sc_hd__inv_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24693_ _25374_/CLK _16104_/X HRESETn VGND VGND VPWR VPWR _24693_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25233__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23644_ _23635_/CLK _19686_/X VGND VGND VPWR VPWR _23644_/Q sky130_fd_sc_hd__dfxtp_4
X_20856_ _24038_/Q VGND VGND VPWR VPWR _20856_/Y sky130_fd_sc_hd__inv_2
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23575_ _23550_/CLK _19881_/X VGND VGND VPWR VPWR _19879_/A sky130_fd_sc_hd__dfxtp_4
X_20787_ _13136_/A _24021_/Q _20783_/B VGND VGND VPWR VPWR _20787_/X sky130_fd_sc_hd__or3_4
XFILLER_23_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25314_ _23904_/CLK _25314_/D HRESETn VGND VGND VPWR VPWR _25314_/Q sky130_fd_sc_hd__dfrtp_4
X_22526_ _22798_/A VGND VGND VPWR VPWR _22526_/X sky130_fd_sc_hd__buf_2
XFILLER_126_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23059__B1 _22798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15536__B2 _15535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25245_ _25070_/CLK _25245_/D HRESETn VGND VGND VPWR VPWR _25245_/Q sky130_fd_sc_hd__dfrtp_4
X_22457_ _20851_/Y _23126_/A _16699_/Y _22271_/X VGND VGND VPWR VPWR _22458_/B sky130_fd_sc_hd__o22a_4
X_12210_ _22400_/A VGND VGND VPWR VPWR _12210_/Y sky130_fd_sc_hd__inv_2
X_21408_ _21408_/A VGND VGND VPWR VPWR _21409_/A sky130_fd_sc_hd__buf_2
X_13190_ _13190_/A _23508_/Q VGND VGND VPWR VPWR _13190_/X sky130_fd_sc_hd__or2_4
X_25176_ _25172_/CLK _14267_/X HRESETn VGND VGND VPWR VPWR _14266_/A sky130_fd_sc_hd__dfrtp_4
X_22388_ _22387_/X VGND VGND VPWR VPWR _22388_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20293__B1 _19995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12770__A1 _25363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12141_ _12128_/B VGND VGND VPWR VPWR _12141_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24127_ _24133_/CLK _18771_/Y HRESETn VGND VGND VPWR VPWR _18688_/A sky130_fd_sc_hd__dfrtp_4
X_21339_ _14428_/Y _21338_/X _14468_/Y _17415_/A VGND VGND VPWR VPWR _21339_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12770__B2 _12769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24186__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12172__C _15652_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22034__A1 _21821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12072_ _16183_/A _12060_/B _12066_/X _12072_/D VGND VGND VPWR VPWR _12072_/X sky130_fd_sc_hd__or4_4
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22034__B2 _22033_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24115__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24058_ _24492_/CLK _20945_/X HRESETn VGND VGND VPWR VPWR _20943_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15900_ _15900_/A VGND VGND VPWR VPWR _15900_/X sky130_fd_sc_hd__buf_2
XANTENNA__22585__A2 _23226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12522__B2 _24858_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23009_ _23009_/A _22394_/X _22812_/C VGND VGND VPWR VPWR _23009_/X sky130_fd_sc_hd__and3_4
X_16880_ _16880_/A VGND VGND VPWR VPWR _16880_/X sky130_fd_sc_hd__buf_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21873__A1_N _12819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15831_ _12324_/Y _15829_/X _15620_/X _15829_/X VGND VGND VPWR VPWR _24814_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15472__B1 _15471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19738__B1 _19715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18550_ _18496_/A _18477_/C VGND VGND VPWR VPWR _18550_/X sky130_fd_sc_hd__or2_4
XFILLER_58_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12974_ _12845_/B _12970_/X VGND VGND VPWR VPWR _12974_/Y sky130_fd_sc_hd__nand2_4
X_15762_ _12514_/Y _15759_/X _15623_/X _15759_/X VGND VGND VPWR VPWR _24848_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17501_ _24299_/Q VGND VGND VPWR VPWR _17630_/A sky130_fd_sc_hd__inv_2
XFILLER_46_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14713_ _14712_/X _13760_/X _14712_/X _13760_/X VGND VGND VPWR VPWR _14713_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11925_ _11924_/X VGND VGND VPWR VPWR _11947_/A sky130_fd_sc_hd__buf_2
X_18481_ _18496_/A _18481_/B _18456_/X _18490_/B VGND VGND VPWR VPWR _18482_/B sky130_fd_sc_hd__or4_4
XFILLER_73_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15693_ _18019_/A VGND VGND VPWR VPWR _15693_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12909__A _12936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17432_ _17432_/A VGND VGND VPWR VPWR _17432_/X sky130_fd_sc_hd__buf_2
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11813__A _11812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11856_ HWDATA[2] VGND VGND VPWR VPWR _11856_/X sky130_fd_sc_hd__buf_2
X_14644_ _13609_/B _14643_/Y _18006_/A _14643_/Y VGND VGND VPWR VPWR _14644_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14575_ _14574_/X _14555_/X _25263_/Q VGND VGND VPWR VPWR _14575_/Y sky130_fd_sc_hd__o21ai_4
X_17363_ _17350_/B _17349_/X _17289_/A _17359_/Y VGND VGND VPWR VPWR _17363_/X sky130_fd_sc_hd__a211o_4
X_11787_ _25525_/Q VGND VGND VPWR VPWR _11787_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19102_ _23845_/Q VGND VGND VPWR VPWR _19102_/Y sky130_fd_sc_hd__inv_2
X_16314_ _16313_/Y _16311_/X _15957_/X _16311_/X VGND VGND VPWR VPWR _24619_/D sky130_fd_sc_hd__a2bb2o_4
X_13526_ _13643_/B VGND VGND VPWR VPWR _13526_/Y sky130_fd_sc_hd__inv_2
X_17294_ _17293_/X VGND VGND VPWR VPWR _17295_/B sky130_fd_sc_hd__inv_2
XFILLER_9_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24956__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19033_ _19032_/Y _19030_/X _18940_/X _19030_/X VGND VGND VPWR VPWR _23870_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21022__A _21015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13457_ _13457_/A _13457_/B _13457_/C VGND VGND VPWR VPWR _13461_/B sky130_fd_sc_hd__and3_4
X_16245_ _16244_/Y _16241_/X _15897_/X _16241_/X VGND VGND VPWR VPWR _24644_/D sky130_fd_sc_hd__a2bb2o_4
X_12408_ _12291_/A _12406_/A VGND VGND VPWR VPWR _12408_/X sky130_fd_sc_hd__or2_4
XFILLER_126_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13388_ _13452_/A _23655_/Q VGND VGND VPWR VPWR _13389_/C sky130_fd_sc_hd__or2_4
X_16176_ _16176_/A VGND VGND VPWR VPWR _16176_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_20_0_HCLK clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_41_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12339_ _12339_/A _12332_/X _12335_/X _12339_/D VGND VGND VPWR VPWR _12339_/X sky130_fd_sc_hd__or4_4
X_15127_ _15422_/A _15125_/Y _24968_/Q _15126_/Y VGND VGND VPWR VPWR _15127_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15955__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16190__A1_N _16189_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15058_ _14986_/A VGND VGND VPWR VPWR _15246_/A sky130_fd_sc_hd__buf_2
X_19935_ _19935_/A VGND VGND VPWR VPWR _19935_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14009_ _14001_/D _14009_/B VGND VGND VPWR VPWR _14010_/C sky130_fd_sc_hd__or2_4
XANTENNA__12513__B2 _24873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19866_ _20338_/A _18278_/D _19888_/C VGND VGND VPWR VPWR _19866_/X sky130_fd_sc_hd__or3_4
XFILLER_64_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20587__A1 _14128_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21784__B1 _13784_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18817_ _18682_/B _18820_/B VGND VGND VPWR VPWR _18817_/Y sky130_fd_sc_hd__nand2_4
X_19797_ _19797_/A VGND VGND VPWR VPWR _19797_/X sky130_fd_sc_hd__buf_2
XANTENNA__16786__A HWDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18748_ _18610_/A _18747_/Y VGND VGND VPWR VPWR _18748_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_144_0_HCLK clkbuf_7_72_0_HCLK/X VGND VGND VPWR VPWR _24209_/CLK sky130_fd_sc_hd__clkbuf_1
X_18679_ _18679_/A VGND VGND VPWR VPWR _18680_/D sky130_fd_sc_hd__inv_2
X_20710_ _22407_/A _20698_/X _20706_/X _20709_/Y VGND VGND VPWR VPWR _20711_/A sky130_fd_sc_hd__o22a_4
XFILLER_24_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21690_ _21539_/X _21592_/X _21646_/X _21689_/X VGND VGND VPWR VPWR HRDATA[2] sky130_fd_sc_hd__or4_4
X_20641_ _20641_/A VGND VGND VPWR VPWR _23976_/D sky130_fd_sc_hd__inv_2
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23360_ _21003_/X VGND VGND VPWR VPWR IRQ[6] sky130_fd_sc_hd__buf_2
X_20572_ _14425_/Y _20556_/X _20546_/X _20571_/X VGND VGND VPWR VPWR _20572_/X sky130_fd_sc_hd__a211o_4
XFILLER_20_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16715__B1 _16442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24697__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22311_ _21826_/A _22311_/B VGND VGND VPWR VPWR _22311_/X sky130_fd_sc_hd__and2_4
XANTENNA__18225__B _18217_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24626__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23291_ _23291_/A _22832_/B VGND VGND VPWR VPWR _23291_/X sky130_fd_sc_hd__or2_4
XANTENNA__16026__A _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25030_ _25029_/CLK _14875_/Y HRESETn VGND VGND VPWR VPWR _14869_/A sky130_fd_sc_hd__dfrtp_4
X_22242_ _22229_/A _20342_/Y VGND VGND VPWR VPWR _22242_/X sky130_fd_sc_hd__or2_4
XANTENNA__12201__B1 _12199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14191__D _13777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22173_ _15465_/Y _21352_/X _14226_/Y _21338_/X VGND VGND VPWR VPWR _22174_/A sky130_fd_sc_hd__o22a_4
XANTENNA__16158__A1_N _16156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21124_ _14492_/Y _21139_/B _14182_/Y _21352_/A VGND VGND VPWR VPWR _21124_/X sky130_fd_sc_hd__o22a_4
XFILLER_99_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13385__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21055_ _21054_/X VGND VGND VPWR VPWR _21055_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20006_ _20006_/A VGND VGND VPWR VPWR _22014_/B sky130_fd_sc_hd__inv_2
XANTENNA__25485__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_40_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_81_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25414__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24814_ _24836_/CLK _24814_/D HRESETn VGND VGND VPWR VPWR _24814_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23306__B _23305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21527__B1 _24809_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21107__A _21069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21957_ _14632_/A _19606_/Y _21958_/A _19604_/Y VGND VGND VPWR VPWR _21957_/X sky130_fd_sc_hd__o22a_4
X_24745_ _24792_/CLK _15976_/X HRESETn VGND VGND VPWR VPWR _22550_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/A VGND VGND VPWR VPWR _16371_/A sky130_fd_sc_hd__buf_2
XANTENNA__18943__B2 _18937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _20882_/X _20907_/Y _24486_/Q _20886_/X VGND VGND VPWR VPWR _20908_/X sky130_fd_sc_hd__a2bb2o_4
X_12690_ _12567_/Y _12674_/B _12648_/A _12688_/B VGND VGND VPWR VPWR _12691_/A sky130_fd_sc_hd__a211o_4
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24676_ _24346_/CLK _24676_/D HRESETn VGND VGND VPWR VPWR _24676_/Q sky130_fd_sc_hd__dfrtp_4
X_21888_ _21887_/X _21888_/B VGND VGND VPWR VPWR _21888_/X sky130_fd_sc_hd__or2_4
XANTENNA__16726__A1_N _15310_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23322__A _22792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23627_ _23635_/CLK _19733_/X VGND VGND VPWR VPWR _23627_/Q sky130_fd_sc_hd__dfxtp_4
X_20839_ _16706_/Y _20836_/X _20824_/X _20838_/X VGND VGND VPWR VPWR _20839_/X sky130_fd_sc_hd__o22a_4
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _14330_/X VGND VGND VPWR VPWR _14360_/X sky130_fd_sc_hd__buf_2
XFILLER_23_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17320__A _17253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23558_ _25246_/CLK _19926_/X VGND VGND VPWR VPWR _19925_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_35_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _13227_/A VGND VGND VPWR VPWR _13312_/A sky130_fd_sc_hd__buf_2
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22509_ _21162_/A _13782_/X _21499_/B VGND VGND VPWR VPWR _22510_/A sky130_fd_sc_hd__or3_4
XFILLER_13_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14291_ _14291_/A _14296_/A _14291_/C _14291_/D VGND VGND VPWR VPWR _14292_/A sky130_fd_sc_hd__or4_4
XFILLER_122_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24367__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23489_ _23609_/CLK _23489_/D VGND VGND VPWR VPWR _23489_/Q sky130_fd_sc_hd__dfxtp_4
X_13242_ _13320_/A _13242_/B VGND VGND VPWR VPWR _13243_/C sky130_fd_sc_hd__or2_4
X_16030_ _16029_/Y _16027_/X _15962_/X _16027_/X VGND VGND VPWR VPWR _24721_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25228_ _23967_/CLK _25228_/D HRESETn VGND VGND VPWR VPWR _13999_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_104_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12743__B2 _24783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13173_ _17453_/A VGND VGND VPWR VPWR _13173_/X sky130_fd_sc_hd__buf_2
X_25159_ _25305_/CLK _14322_/X HRESETn VGND VGND VPWR VPWR _25159_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12124_ _12123_/Y _12119_/X _11867_/X _12119_/X VGND VGND VPWR VPWR _12124_/X sky130_fd_sc_hd__a2bb2o_4
X_17981_ _18087_/A VGND VGND VPWR VPWR _18201_/A sky130_fd_sc_hd__buf_2
XFILLER_105_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19720_ _19706_/Y VGND VGND VPWR VPWR _19720_/X sky130_fd_sc_hd__buf_2
X_12055_ _12054_/X VGND VGND VPWR VPWR _12060_/B sky130_fd_sc_hd__buf_2
X_16932_ _16925_/X _16932_/B _16930_/X _16932_/D VGND VGND VPWR VPWR _16932_/X sky130_fd_sc_hd__or4_4
XANTENNA__17990__A _17990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11808__A HWDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19651_ _19650_/Y _19646_/X _19599_/X _19646_/X VGND VGND VPWR VPWR _23656_/D sky130_fd_sc_hd__a2bb2o_4
X_16863_ _19777_/A VGND VGND VPWR VPWR _16863_/X sky130_fd_sc_hd__buf_2
XANTENNA__23931__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18602_ _16608_/A _18782_/A _16555_/Y _18719_/A VGND VGND VPWR VPWR _18602_/X sky130_fd_sc_hd__a2bb2o_4
X_15814_ _12337_/Y _15812_/X _11788_/X _15812_/X VGND VGND VPWR VPWR _24825_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19582_ _13815_/A _21143_/A VGND VGND VPWR VPWR _19582_/X sky130_fd_sc_hd__or2_4
XFILLER_111_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16794_ _24432_/Q VGND VGND VPWR VPWR _16794_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23216__B _21519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18533_ _18420_/Y _18540_/A _18461_/Y _18542_/B VGND VGND VPWR VPWR _18539_/B sky130_fd_sc_hd__or4_4
XANTENNA__21017__A _25355_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15745_ HWDATA[14] VGND VGND VPWR VPWR _15745_/X sky130_fd_sc_hd__buf_2
XFILLER_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12957_ _12944_/B _12944_/D _12884_/A _12953_/Y VGND VGND VPWR VPWR _12957_/X sky130_fd_sc_hd__a211o_4
XFILLER_34_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12639__A _12631_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_217_0_HCLK clkbuf_8_217_0_HCLK/A VGND VGND VPWR VPWR _24413_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_34_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22730__A2 _22419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11908_ _13678_/B _11879_/B _11896_/X _11871_/A VGND VGND VPWR VPWR _11908_/X sky130_fd_sc_hd__a211o_4
X_18464_ _18405_/Y _18461_/Y _18464_/C _18464_/D VGND VGND VPWR VPWR _18465_/C sky130_fd_sc_hd__or4_4
X_15676_ _15643_/Y _15669_/X _15647_/X _24877_/Q _15675_/X VGND VGND VPWR VPWR _24877_/D
+ sky130_fd_sc_hd__a32o_4
X_12888_ _12841_/B _12887_/X VGND VGND VPWR VPWR _12889_/A sky130_fd_sc_hd__or2_4
X_17415_ _17415_/A VGND VGND VPWR VPWR _17416_/A sky130_fd_sc_hd__buf_2
XANTENNA__23232__A _23232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14627_ _21962_/A _13638_/X _14626_/A _13637_/A VGND VGND VPWR VPWR _14628_/A sky130_fd_sc_hd__o22a_4
X_11839_ _11835_/Y _11836_/X _11838_/X _11836_/X VGND VGND VPWR VPWR _11839_/X sky130_fd_sc_hd__a2bb2o_4
X_18395_ _16202_/Y _18459_/A _16202_/Y _18459_/A VGND VGND VPWR VPWR _18395_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17346_ _17243_/D _17346_/B VGND VGND VPWR VPWR _17347_/B sky130_fd_sc_hd__or2_4
X_14558_ _14558_/A VGND VGND VPWR VPWR _14558_/X sky130_fd_sc_hd__buf_2
XFILLER_18_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24790__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18162__A2 _18146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13509_ _13509_/A VGND VGND VPWR VPWR _13509_/Y sky130_fd_sc_hd__inv_2
X_17277_ _17194_/Y _17277_/B VGND VGND VPWR VPWR _17278_/C sky130_fd_sc_hd__or2_4
X_14489_ _14487_/Y _14488_/X _14395_/X _14488_/X VGND VGND VPWR VPWR _25103_/D sky130_fd_sc_hd__a2bb2o_4
X_19016_ _19030_/A VGND VGND VPWR VPWR _19016_/X sky130_fd_sc_hd__buf_2
X_16228_ _11800_/A VGND VGND VPWR VPWR _16228_/X sky130_fd_sc_hd__buf_2
XANTENNA__24037__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13189__B _23908_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16159_ _21691_/A VGND VGND VPWR VPWR _16159_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18996__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19918_ _19918_/A VGND VGND VPWR VPWR _19918_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19849_ _23587_/Q VGND VGND VPWR VPWR _19849_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21221__A2 _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21703__A1_N _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_27_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22860_ _22860_/A _22626_/B VGND VGND VPWR VPWR _22860_/X sky130_fd_sc_hd__or2_4
X_21811_ _21648_/A _21811_/B VGND VGND VPWR VPWR _21811_/X sky130_fd_sc_hd__or2_4
X_22791_ _20749_/Y _22280_/X _20888_/Y _22790_/X VGND VGND VPWR VPWR _22791_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12549__A _24851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24530_ _24553_/CLK _24530_/D HRESETn VGND VGND VPWR VPWR _24530_/Q sky130_fd_sc_hd__dfrtp_4
X_21742_ _20828_/Y _21588_/X _24000_/Q _21589_/X VGND VGND VPWR VPWR _21742_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24878__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12239__A2_N _24749_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24461_ _24462_/CLK _24461_/D HRESETn VGND VGND VPWR VPWR _24461_/Q sky130_fd_sc_hd__dfrtp_4
X_21673_ _21449_/A _19482_/Y VGND VGND VPWR VPWR _21675_/B sky130_fd_sc_hd__or2_4
XANTENNA__24807__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23412_ _23533_/CLK _23412_/D VGND VGND VPWR VPWR _20315_/A sky130_fd_sc_hd__dfxtp_4
X_20624_ _23973_/Q _20621_/A VGND VGND VPWR VPWR _20624_/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24392_ _24806_/CLK _24392_/D HRESETn VGND VGND VPWR VPWR _21004_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_123_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23343_ _23343_/A _23343_/B VGND VGND VPWR VPWR _23343_/X sky130_fd_sc_hd__and2_4
X_20555_ _20554_/X VGND VGND VPWR VPWR _23935_/D sky130_fd_sc_hd__inv_2
XANTENNA__24460__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23274_ _23274_/A _23274_/B VGND VGND VPWR VPWR _23281_/C sky130_fd_sc_hd__and2_4
X_20486_ _20479_/A _20486_/B _24070_/Q VGND VGND VPWR VPWR _20486_/X sky130_fd_sc_hd__and3_4
XANTENNA__20248__B1 _18267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25013_ _25016_/CLK _15225_/X HRESETn VGND VGND VPWR VPWR _25013_/Q sky130_fd_sc_hd__dfrtp_4
X_22225_ _21192_/A VGND VGND VPWR VPWR _22229_/A sky130_fd_sc_hd__buf_2
XFILLER_69_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22156_ _16608_/A _21323_/X _15667_/A _22155_/X VGND VGND VPWR VPWR _22157_/C sky130_fd_sc_hd__a211o_4
XANTENNA__18861__B1 _16457_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_109_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_219_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21107_ _21069_/A VGND VGND VPWR VPWR _21108_/B sky130_fd_sc_hd__buf_2
XFILLER_105_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22087_ _23085_/A _22087_/B _22086_/X VGND VGND VPWR VPWR _22087_/X sky130_fd_sc_hd__and3_4
XFILLER_121_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12489__B1 _12394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21038_ _21006_/A _21038_/B VGND VGND VPWR VPWR _21038_/X sky130_fd_sc_hd__and2_4
XANTENNA__18613__B1 _24529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13860_ _23990_/Q VGND VGND VPWR VPWR _13860_/X sky130_fd_sc_hd__buf_2
XFILLER_74_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12811_ _12850_/B _12792_/A _25376_/Q _12758_/Y VGND VGND VPWR VPWR _12815_/C sky130_fd_sc_hd__a2bb2o_4
X_13791_ _13815_/A _14255_/A VGND VGND VPWR VPWR _13791_/X sky130_fd_sc_hd__or2_4
XANTENNA__23224__A1_N _17261_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22989_ _20771_/Y _22988_/X _20910_/Y _21211_/X VGND VGND VPWR VPWR _22990_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22173__B1 _14226_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21515__A3 _21514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15530_ _15528_/Y _15524_/X HADDR[7] _15529_/X VGND VGND VPWR VPWR _15530_/X sky130_fd_sc_hd__a2bb2o_4
X_12742_ _25366_/Q VGND VGND VPWR VPWR _12842_/A sky130_fd_sc_hd__inv_2
X_24728_ _24345_/CLK _16013_/X HRESETn VGND VGND VPWR VPWR _16012_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_190_0_HCLK clkbuf_7_95_0_HCLK/X VGND VGND VPWR VPWR _25433_/CLK sky130_fd_sc_hd__clkbuf_1
X_12673_ _12672_/X VGND VGND VPWR VPWR _25408_/D sky130_fd_sc_hd__inv_2
X_15461_ _24945_/Q VGND VGND VPWR VPWR _15461_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12609__D _12567_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24548__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24659_ _24654_/CLK _24659_/D HRESETn VGND VGND VPWR VPWR _23129_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18146__A _17928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _21531_/A _17199_/A _16361_/Y _17199_/Y VGND VGND VPWR VPWR _17201_/D sky130_fd_sc_hd__o22a_4
XFILLER_54_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_47_0_HCLK clkbuf_8_47_0_HCLK/A VGND VGND VPWR VPWR _23384_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _14405_/Y _14409_/X _14411_/X _14409_/X VGND VGND VPWR VPWR _25132_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _18180_/A _23862_/Q VGND VGND VPWR VPWR _18181_/C sky130_fd_sc_hd__or2_4
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ _15392_/A _15408_/A VGND VGND VPWR VPWR _15392_/X sky130_fd_sc_hd__or2_4
XFILLER_15_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17131_ _16960_/Y _17151_/A VGND VGND VPWR VPWR _17148_/A sky130_fd_sc_hd__or2_4
XFILLER_11_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14343_ _14339_/Y _14336_/C VGND VGND VPWR VPWR _14348_/A sky130_fd_sc_hd__or2_4
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14274_ _14273_/Y _14271_/X _14239_/X _14271_/X VGND VGND VPWR VPWR _14274_/X sky130_fd_sc_hd__a2bb2o_4
X_17062_ _16981_/A _17061_/Y VGND VGND VPWR VPWR _17062_/X sky130_fd_sc_hd__or2_4
XANTENNA__24130__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20239__B1 _19758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13225_ _13225_/A VGND VGND VPWR VPWR _13310_/A sky130_fd_sc_hd__buf_2
X_16013_ _16012_/Y _16010_/X _11764_/X _16010_/X VGND VGND VPWR VPWR _16013_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13156_ _13155_/Y VGND VGND VPWR VPWR _13156_/X sky130_fd_sc_hd__buf_2
XFILLER_48_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14943__A2_N _14941_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12107_ _12119_/A VGND VGND VPWR VPWR _12107_/X sky130_fd_sc_hd__buf_2
XANTENNA__25336__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13087_ _12992_/Y _13086_/X VGND VGND VPWR VPWR _13087_/X sky130_fd_sc_hd__or2_4
X_17964_ _14785_/A VGND VGND VPWR VPWR _18217_/A sky130_fd_sc_hd__buf_2
XFILLER_97_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19703_ _19702_/Y _19697_/X _19658_/X _19697_/A VGND VGND VPWR VPWR _23637_/D sky130_fd_sc_hd__a2bb2o_4
X_12038_ _25478_/Q VGND VGND VPWR VPWR _12038_/Y sky130_fd_sc_hd__inv_2
X_16915_ _22902_/A _24264_/Q _16117_/Y _16914_/Y VGND VGND VPWR VPWR _16922_/A sky130_fd_sc_hd__o22a_4
XANTENNA__18604__B1 _16560_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17895_ _17909_/A _17894_/X VGND VGND VPWR VPWR _17895_/Y sky130_fd_sc_hd__nand2_4
XFILLER_66_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19634_ _23661_/Q VGND VGND VPWR VPWR _21177_/B sky130_fd_sc_hd__inv_2
XFILLER_65_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22951__A2 _22833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16846_ _14945_/Y _16844_/X _16528_/X _16844_/X VGND VGND VPWR VPWR _16846_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16091__B1 _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19565_ _22229_/B _19562_/X _11934_/X _19562_/X VGND VGND VPWR VPWR _19565_/X sky130_fd_sc_hd__a2bb2o_4
X_16777_ _16776_/Y _16773_/X _16521_/X _16773_/X VGND VGND VPWR VPWR _16777_/X sky130_fd_sc_hd__a2bb2o_4
X_13989_ _13989_/A VGND VGND VPWR VPWR _13989_/X sky130_fd_sc_hd__buf_2
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18516_ _24168_/Q _18519_/B VGND VGND VPWR VPWR _18516_/X sky130_fd_sc_hd__or2_4
X_15728_ _15728_/A VGND VGND VPWR VPWR _15728_/X sky130_fd_sc_hd__buf_2
X_19496_ _22325_/B _19495_/X _11930_/X _19495_/X VGND VGND VPWR VPWR _23708_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24971__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21911__B1 _21270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18447_ _23232_/A _18456_/A _16258_/Y _24149_/Q VGND VGND VPWR VPWR _18447_/X sky130_fd_sc_hd__a2bb2o_4
X_15659_ _16640_/B _15777_/B VGND VGND VPWR VPWR _15659_/X sky130_fd_sc_hd__or2_4
XANTENNA__24289__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24900__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18378_ _18376_/Y _18372_/X _24182_/Q _18377_/X VGND VGND VPWR VPWR _18378_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17329_ _17252_/B _17307_/X VGND VGND VPWR VPWR _17330_/A sky130_fd_sc_hd__or2_4
XANTENNA__11720__B _11720_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14157__B1 _25123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20340_ _20339_/Y VGND VGND VPWR VPWR _20340_/X sky130_fd_sc_hd__buf_2
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20271_ _21252_/B _20266_/X _19841_/A _20266_/A VGND VGND VPWR VPWR _23429_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22010_ _22024_/A _22010_/B VGND VGND VPWR VPWR _22010_/X sky130_fd_sc_hd__or2_4
XFILLER_118_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25077__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25006__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23961_ _24955_/CLK _21001_/X HRESETn VGND VGND VPWR VPWR _14249_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22912_ _22907_/X _22910_/X _23117_/C VGND VGND VPWR VPWR _22912_/X sky130_fd_sc_hd__or3_4
X_23892_ _23869_/CLK _18968_/X VGND VGND VPWR VPWR _23892_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22843_ _21530_/X VGND VGND VPWR VPWR _22843_/X sky130_fd_sc_hd__buf_2
XANTENNA__22155__B1 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12178__A2_N _24746_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22695__B _22695_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22774_ _22774_/A _22644_/B VGND VGND VPWR VPWR _22774_/X sky130_fd_sc_hd__or2_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_200_0_HCLK clkbuf_8_201_0_HCLK/A VGND VGND VPWR VPWR _24699_/CLK sky130_fd_sc_hd__clkbuf_1
X_21725_ _18381_/Y _12072_/D _12116_/Y _21561_/X VGND VGND VPWR VPWR _21725_/X sky130_fd_sc_hd__o22a_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24513_ _24545_/CLK _16596_/X HRESETn VGND VGND VPWR VPWR _16594_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24641__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25493_ _24923_/CLK _25493_/D HRESETn VGND VGND VPWR VPWR _11941_/A sky130_fd_sc_hd__dfrtp_4
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_6_0_HCLK clkbuf_8_7_0_HCLK/A VGND VGND VPWR VPWR _23453_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21656_ _21460_/A _21654_/X _21656_/C VGND VGND VPWR VPWR _21656_/X sky130_fd_sc_hd__and3_4
X_24444_ _25002_/CLK _16771_/X HRESETn VGND VGND VPWR VPWR _24444_/Q sky130_fd_sc_hd__dfrtp_4
X_20607_ _14868_/Y _20605_/X _20662_/A _20606_/X VGND VGND VPWR VPWR _20607_/X sky130_fd_sc_hd__a211o_4
XFILLER_21_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24375_ _24376_/CLK _24375_/D HRESETn VGND VGND VPWR VPWR _17031_/A sky130_fd_sc_hd__dfrtp_4
X_21587_ _21408_/A VGND VGND VPWR VPWR _21587_/X sky130_fd_sc_hd__buf_2
XANTENNA__17334__B1 _17279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23326_ _22701_/A _23323_/X _23326_/C VGND VGND VPWR VPWR _23331_/C sky130_fd_sc_hd__and3_4
X_20538_ _20562_/A VGND VGND VPWR VPWR _20558_/C sky130_fd_sc_hd__buf_2
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23257_ _15005_/A _23019_/B _23019_/C VGND VGND VPWR VPWR _23257_/X sky130_fd_sc_hd__and3_4
X_20469_ _20469_/A _24073_/Q VGND VGND VPWR VPWR _20469_/X sky130_fd_sc_hd__or2_4
X_13010_ _13010_/A _13004_/B _13009_/X VGND VGND VPWR VPWR _13011_/A sky130_fd_sc_hd__or3_4
X_22208_ _21595_/A _22208_/B VGND VGND VPWR VPWR _22208_/X sky130_fd_sc_hd__or2_4
XANTENNA__22630__B2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23188_ _22975_/X _23187_/X _23044_/X _11756_/A _23111_/X VGND VGND VPWR VPWR _23188_/X
+ sky130_fd_sc_hd__a32o_4
X_22139_ _15708_/A _22137_/X _22466_/A VGND VGND VPWR VPWR _22139_/X sky130_fd_sc_hd__and3_4
XFILLER_79_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14961_ _14960_/Y VGND VGND VPWR VPWR _14961_/X sky130_fd_sc_hd__buf_2
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16700_ _16645_/A VGND VGND VPWR VPWR _16700_/X sky130_fd_sc_hd__buf_2
X_13912_ _13918_/A _13898_/Y _13908_/X _13918_/C _13911_/X VGND VGND VPWR VPWR _13912_/X
+ sky130_fd_sc_hd__a32o_4
X_17680_ _17494_/Y _17685_/A VGND VGND VPWR VPWR _17682_/B sky130_fd_sc_hd__nand2_4
X_14892_ _25001_/Q _14890_/Y _15187_/A _14905_/A VGND VGND VPWR VPWR _14892_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16631_ _16629_/Y _16630_/Y _16634_/B VGND VGND VPWR VPWR _16631_/X sky130_fd_sc_hd__or3_4
XFILLER_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_10_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_13843_ _13821_/A VGND VGND VPWR VPWR _13843_/X sky130_fd_sc_hd__buf_2
XFILLER_35_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24729__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15820__B1 _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19350_ _19348_/Y _19346_/X _19349_/X _19346_/X VGND VGND VPWR VPWR _19350_/X sky130_fd_sc_hd__a2bb2o_4
X_16562_ _24526_/Q VGND VGND VPWR VPWR _16562_/Y sky130_fd_sc_hd__inv_2
X_13774_ _13593_/X VGND VGND VPWR VPWR _13774_/Y sky130_fd_sc_hd__inv_2
X_18301_ _18303_/B _18301_/B VGND VGND VPWR VPWR _18301_/X sky130_fd_sc_hd__and2_4
X_15513_ _11728_/A VGND VGND VPWR VPWR _15513_/Y sky130_fd_sc_hd__inv_2
X_12725_ _12704_/X _12725_/B _12721_/X VGND VGND VPWR VPWR _25393_/D sky130_fd_sc_hd__and3_4
X_19281_ _21381_/B _19278_/X _16888_/X _19278_/X VGND VGND VPWR VPWR _19281_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16493_ _24552_/Q VGND VGND VPWR VPWR _16493_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24382__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18232_ _18249_/A VGND VGND VPWR VPWR _18233_/A sky130_fd_sc_hd__buf_2
XANTENNA__14387__B1 _13837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11821__A HWDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15444_ _15452_/A VGND VGND VPWR VPWR _15444_/X sky130_fd_sc_hd__buf_2
X_12656_ _12656_/A _12656_/B VGND VGND VPWR VPWR _12656_/Y sky130_fd_sc_hd__nand2_4
XFILLER_129_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12937__A1 _12799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18163_ _17963_/X _18162_/X _24231_/Q _18021_/X VGND VGND VPWR VPWR _24231_/D sky130_fd_sc_hd__o22a_4
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12587_ _25408_/Q VGND VGND VPWR VPWR _12611_/B sky130_fd_sc_hd__inv_2
X_15375_ _15372_/A _15365_/B _15375_/C VGND VGND VPWR VPWR _24978_/D sky130_fd_sc_hd__and3_4
XFILLER_15_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17114_ _17031_/A _17114_/B VGND VGND VPWR VPWR _17115_/C sky130_fd_sc_hd__or2_4
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14326_ _25156_/Q _12163_/X _14325_/X VGND VGND VPWR VPWR _14327_/A sky130_fd_sc_hd__a21o_4
X_18094_ _18056_/A _18094_/B VGND VGND VPWR VPWR _18094_/X sky130_fd_sc_hd__or2_4
X_17045_ _17045_/A _17041_/X _17045_/C VGND VGND VPWR VPWR _17045_/X sky130_fd_sc_hd__or3_4
XANTENNA__19078__B1 _19077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25517__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14257_ _14257_/A VGND VGND VPWR VPWR _14258_/A sky130_fd_sc_hd__buf_2
X_13208_ _13155_/Y VGND VGND VPWR VPWR _13457_/A sky130_fd_sc_hd__buf_2
XANTENNA__18825__B1 _16501_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14188_ _12052_/A _15549_/B VGND VGND VPWR VPWR _16369_/D sky130_fd_sc_hd__or2_4
XFILLER_48_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15639__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23116__A1_N _17239_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13139_ _20675_/B VGND VGND VPWR VPWR _13139_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18996_ HWDATA[5] VGND VGND VPWR VPWR _18996_/X sky130_fd_sc_hd__buf_2
X_17947_ _17957_/A _17945_/X _17947_/C VGND VGND VPWR VPWR _17947_/X sky130_fd_sc_hd__and3_4
XFILLER_26_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17878_ _16920_/Y _17878_/B VGND VGND VPWR VPWR _17878_/X sky130_fd_sc_hd__or2_4
XFILLER_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16829_ _24415_/Q VGND VGND VPWR VPWR _16829_/Y sky130_fd_sc_hd__inv_2
X_19617_ _19617_/A VGND VGND VPWR VPWR _19617_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12099__A _16183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15811__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19548_ _19546_/Y _19544_/X _19547_/X _19544_/X VGND VGND VPWR VPWR _23689_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25288__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19479_ _21941_/B _19476_/X _11943_/X _19476_/X VGND VGND VPWR VPWR _23713_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21510_ _21510_/A _21407_/X _21510_/C _21509_/X VGND VGND VPWR VPWR HRDATA[1] sky130_fd_sc_hd__or4_4
X_22490_ _12220_/X _22489_/X _16918_/A _21045_/X VGND VGND VPWR VPWR _22490_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24052__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_30_0_HCLK clkbuf_8_31_0_HCLK/A VGND VGND VPWR VPWR _24373_/CLK sky130_fd_sc_hd__clkbuf_1
X_21441_ _16927_/X _22821_/A _12280_/Y _22429_/A VGND VGND VPWR VPWR _21441_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21859__B _21859_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_93_0_HCLK clkbuf_8_93_0_HCLK/A VGND VGND VPWR VPWR _24136_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24160_ _24541_/CLK _18546_/X HRESETn VGND VGND VPWR VPWR _24160_/Q sky130_fd_sc_hd__dfrtp_4
X_21372_ _21372_/A VGND VGND VPWR VPWR _21393_/A sky130_fd_sc_hd__buf_2
XANTENNA__15878__B1 _11774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23111_ _15544_/X VGND VGND VPWR VPWR _23111_/X sky130_fd_sc_hd__buf_2
X_20323_ _20317_/X _19586_/D _11838_/A _21978_/B _20326_/A VGND VGND VPWR VPWR _20323_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25258__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19069__B1 _18997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24091_ _25246_/CLK _20959_/X HRESETn VGND VGND VPWR VPWR _12019_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16034__A _15995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23042_ _23041_/X VGND VGND VPWR VPWR _23042_/Y sky130_fd_sc_hd__inv_2
X_20254_ _20266_/A VGND VGND VPWR VPWR _20254_/X sky130_fd_sc_hd__buf_2
XANTENNA__15893__A3 _11812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12281__B _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20185_ _20184_/Y _20182_/X _20099_/X _20182_/X VGND VGND VPWR VPWR _20185_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24993_ _24984_/CLK _24993_/D HRESETn VGND VGND VPWR VPWR _15155_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13393__A _13457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23944_ _25205_/CLK _23944_/D HRESETn VGND VGND VPWR VPWR _18884_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24893__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16055__B1 _15758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24822__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23875_ _25485_/CLK _23875_/D VGND VGND VPWR VPWR _19020_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_71_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23314__B _23314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22826_ _23069_/B VGND VGND VPWR VPWR _22826_/X sky130_fd_sc_hd__buf_2
XFILLER_60_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22757_ _22756_/X VGND VGND VPWR VPWR _22758_/D sky130_fd_sc_hd__inv_2
XANTENNA__16341__A2_N _16337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16209__A _23004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12510_ _12510_/A VGND VGND VPWR VPWR _12510_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15719__A1_N _12546_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13490_ _13488_/Y _13489_/X _11858_/X _13489_/X VGND VGND VPWR VPWR _25306_/D sky130_fd_sc_hd__a2bb2o_4
X_21708_ _21708_/A _14258_/A VGND VGND VPWR VPWR _21712_/A sky130_fd_sc_hd__or2_4
XFILLER_40_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25476_ _25461_/CLK _25476_/D HRESETn VGND VGND VPWR VPWR _25476_/Q sky130_fd_sc_hd__dfrtp_4
X_22688_ _13562_/Y _22726_/B VGND VGND VPWR VPWR _22688_/X sky130_fd_sc_hd__and2_4
X_12441_ _12286_/C _12440_/X _12394_/X VGND VGND VPWR VPWR _12441_/Y sky130_fd_sc_hd__a21oi_4
X_21639_ _23671_/Q _21362_/X _23687_/Q _22390_/B VGND VGND VPWR VPWR _21639_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24427_ _24427_/CLK _24427_/D HRESETn VGND VGND VPWR VPWR _24427_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18646__A1_N _16590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12372_ _25325_/Q VGND VGND VPWR VPWR _12378_/A sky130_fd_sc_hd__inv_2
X_15160_ _15406_/A _15077_/A _15159_/X _24570_/Q VGND VGND VPWR VPWR _15160_/X sky130_fd_sc_hd__a2bb2o_4
X_24358_ _24612_/CLK _24358_/D HRESETn VGND VGND VPWR VPWR _24358_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_5_1_0_HCLK clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_14111_ _14108_/X VGND VGND VPWR VPWR _14111_/X sky130_fd_sc_hd__buf_2
X_15091_ _24984_/Q _15089_/Y _24990_/Q _15090_/Y VGND VGND VPWR VPWR _15091_/X sky130_fd_sc_hd__a2bb2o_4
X_23309_ _23308_/X VGND VGND VPWR VPWR _23309_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15333__A2 _15316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12472__A _12220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24289_ _24278_/CLK _17671_/X HRESETn VGND VGND VPWR VPWR _24289_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14042_ _14042_/A _14006_/B _25221_/Q _14042_/D VGND VGND VPWR VPWR _14043_/A sky130_fd_sc_hd__or4_4
XFILLER_69_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22603__A1 _17744_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22603__B2 _22429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18850_ _16481_/Y _18647_/X _16481_/Y _18647_/X VGND VGND VPWR VPWR _18854_/A sky130_fd_sc_hd__a2bb2o_4
X_17801_ _17792_/X VGND VGND VPWR VPWR _17805_/B sky130_fd_sc_hd__inv_2
XFILLER_95_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16294__B1 _15944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18781_ _18619_/Y VGND VGND VPWR VPWR _18792_/B sky130_fd_sc_hd__buf_2
X_15993_ _16276_/B VGND VGND VPWR VPWR _15993_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23208__C _23203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17732_ _21491_/A _17731_/X _21491_/A _17731_/X VGND VGND VPWR VPWR _17733_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14944_ _14944_/A VGND VGND VPWR VPWR _14944_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20917__B2 _20913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17663_ _17576_/Y _17662_/X VGND VGND VPWR VPWR _17683_/A sky130_fd_sc_hd__or2_4
X_14875_ _14874_/X VGND VGND VPWR VPWR _14875_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22119__B1 _22087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24563__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19402_ _19398_/Y _19401_/X _19313_/X _19401_/X VGND VGND VPWR VPWR _23740_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21590__B2 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16614_ _16550_/A VGND VGND VPWR VPWR _16614_/X sky130_fd_sc_hd__buf_2
XFILLER_1_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13826_ _13569_/Y _13822_/X _11809_/X _13825_/X VGND VGND VPWR VPWR _13826_/X sky130_fd_sc_hd__a2bb2o_4
X_17594_ _17584_/C _17604_/A VGND VGND VPWR VPWR _17597_/B sky130_fd_sc_hd__or2_4
XFILLER_90_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19333_ _19332_/X VGND VGND VPWR VPWR _19333_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16545_ _16545_/A VGND VGND VPWR VPWR _16545_/X sky130_fd_sc_hd__buf_2
X_13757_ _13757_/A _13757_/B VGND VGND VPWR VPWR _13758_/B sky130_fd_sc_hd__and2_4
XANTENNA__17546__B1 _11860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15023__A _15023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12708_ _12708_/A _12708_/B VGND VGND VPWR VPWR _12712_/B sky130_fd_sc_hd__or2_4
X_19264_ _13736_/X _19084_/D _19845_/C VGND VGND VPWR VPWR _19264_/X sky130_fd_sc_hd__or3_4
X_16476_ _16476_/A VGND VGND VPWR VPWR _16476_/Y sky130_fd_sc_hd__inv_2
X_13688_ _11685_/Y _13688_/B VGND VGND VPWR VPWR _13689_/B sky130_fd_sc_hd__or2_4
XANTENNA__12180__A1_N _12179_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18215_ _18215_/A _19009_/A VGND VGND VPWR VPWR _18216_/C sky130_fd_sc_hd__or2_4
X_15427_ _15426_/X VGND VGND VPWR VPWR _15427_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_17_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_34_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_12639_ _12631_/B VGND VGND VPWR VPWR _12648_/A sky130_fd_sc_hd__buf_2
X_19195_ _19195_/A VGND VGND VPWR VPWR _19195_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13032__B1 _13031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18146_ _17928_/A _18146_/B _18146_/C VGND VGND VPWR VPWR _18146_/X sky130_fd_sc_hd__and3_4
X_15358_ _15298_/B _15352_/X _15318_/A _15355_/B VGND VGND VPWR VPWR _15359_/A sky130_fd_sc_hd__a211o_4
XFILLER_116_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14309_ _14306_/X _14308_/Y _25311_/Q _14306_/X VGND VGND VPWR VPWR _25165_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25351__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18077_ _18224_/A _18072_/X _18077_/C VGND VGND VPWR VPWR _18078_/C sky130_fd_sc_hd__or3_4
XFILLER_85_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15289_ _15285_/X VGND VGND VPWR VPWR _15346_/A sky130_fd_sc_hd__buf_2
X_17028_ _24385_/Q VGND VGND VPWR VPWR _17029_/A sky130_fd_sc_hd__inv_2
XANTENNA__15875__A3 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18979_ _18976_/Y _18972_/X _18977_/X _18978_/X VGND VGND VPWR VPWR _18979_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11726__A _24919_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19223__B1 _19155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21990_ _17900_/A _20331_/A _17887_/Y _21977_/B VGND VGND VPWR VPWR _21990_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20908__B2 _20886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20941_ _20818_/X _20940_/Y _24494_/Q _20864_/X VGND VGND VPWR VPWR _20941_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17413__A _17413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20872_ _20860_/X _20871_/Y _24478_/Q _20865_/X VGND VGND VPWR VPWR _24041_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_82_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24233__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23660_ _23660_/CLK _23660_/D VGND VGND VPWR VPWR _13159_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22611_ _22574_/A _22608_/X _22611_/C VGND VGND VPWR VPWR _22611_/X sky130_fd_sc_hd__and3_4
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23591_ _24089_/CLK _23591_/D VGND VGND VPWR VPWR _19835_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16029__A _16029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22542_ _16597_/A _23226_/B _21731_/X _22541_/X VGND VGND VPWR VPWR _22543_/C sky130_fd_sc_hd__a211o_4
XFILLER_35_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25330_ _25330_/CLK _13095_/X HRESETn VGND VGND VPWR VPWR _25330_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23150__A _22186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22473_ _22470_/X _22472_/X _21416_/X _24851_/Q _22540_/A VGND VGND VPWR VPWR _22473_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25439__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25261_ _25246_/CLK _25261_/D HRESETn VGND VGND VPWR VPWR _13799_/A sky130_fd_sc_hd__dfrtp_4
X_21424_ _21071_/A VGND VGND VPWR VPWR _21525_/A sky130_fd_sc_hd__buf_2
X_24212_ _25508_/CLK _18263_/X HRESETn VGND VGND VPWR VPWR _18259_/A sky130_fd_sc_hd__dfrtp_4
X_25192_ _25192_/CLK _14211_/X HRESETn VGND VGND VPWR VPWR _14209_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25092__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24143_ _24133_/CLK _18709_/Y HRESETn VGND VGND VPWR VPWR _18671_/A sky130_fd_sc_hd__dfrtp_4
X_21355_ _21355_/A VGND VGND VPWR VPWR _21549_/B sky130_fd_sc_hd__buf_2
XFILLER_107_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20306_ _23416_/Q VGND VGND VPWR VPWR _21935_/B sky130_fd_sc_hd__inv_2
XANTENNA__25021__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15866__A3 _15714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24074_ _24069_/CLK _24074_/D HRESETn VGND VGND VPWR VPWR _20469_/A sky130_fd_sc_hd__dfrtp_4
X_21286_ _21278_/X _21286_/B _21290_/C VGND VGND VPWR VPWR _21286_/X sky130_fd_sc_hd__and3_4
XFILLER_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23025_ _12824_/Y _22707_/X _22272_/X _12586_/Y _22844_/X VGND VGND VPWR VPWR _23025_/X
+ sky130_fd_sc_hd__o32a_4
X_20237_ _13266_/B VGND VGND VPWR VPWR _20237_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20168_ _20043_/C _13752_/X _20043_/A _13762_/A VGND VGND VPWR VPWR _20169_/A sky130_fd_sc_hd__or4_4
XANTENNA__17307__B _17249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20014__A _20014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23010__A1 _24725_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12990_ _13048_/A _12990_/B _12990_/C VGND VGND VPWR VPWR _13028_/D sky130_fd_sc_hd__or3_4
X_20099_ _20099_/A VGND VGND VPWR VPWR _20099_/X sky130_fd_sc_hd__buf_2
X_24976_ _24977_/CLK _24976_/D HRESETn VGND VGND VPWR VPWR _15382_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16028__B1 _15959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11941_ _11941_/A VGND VGND VPWR VPWR _11948_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23927_ _25199_/CLK _20973_/X HRESETn VGND VGND VPWR VPWR _20977_/B sky130_fd_sc_hd__dfstp_4
XFILLER_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14660_ _13624_/A VGND VGND VPWR VPWR _19014_/B sky130_fd_sc_hd__buf_2
X_11872_ _11871_/Y VGND VGND VPWR VPWR _11872_/X sky130_fd_sc_hd__buf_2
X_23858_ _23441_/CLK _23858_/D VGND VGND VPWR VPWR _19067_/A sky130_fd_sc_hd__dfxtp_4
X_13611_ _18088_/A VGND VGND VPWR VPWR _17929_/A sky130_fd_sc_hd__buf_2
XANTENNA__19517__B2 _19516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22809_ _22809_/A _22722_/B VGND VGND VPWR VPWR _22814_/B sky130_fd_sc_hd__or2_4
X_14591_ _14571_/Y _14586_/X _14589_/X _14590_/X _14570_/A VGND VGND VPWR VPWR _25080_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_60_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23789_ _23846_/CLK _19261_/X VGND VGND VPWR VPWR _19260_/A sky130_fd_sc_hd__dfxtp_4
X_16330_ _16324_/A VGND VGND VPWR VPWR _16330_/X sky130_fd_sc_hd__buf_2
XFILLER_125_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13542_ _17911_/A _13541_/X VGND VGND VPWR VPWR _13590_/A sky130_fd_sc_hd__and2_4
XFILLER_125_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25528_ _25436_/CLK _25528_/D HRESETn VGND VGND VPWR VPWR _11776_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23956__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16261_ _24637_/Q VGND VGND VPWR VPWR _16261_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23077__A1 _12277_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13473_ _13465_/Y _13471_/Y _13472_/X _13471_/Y VGND VGND VPWR VPWR _13473_/X sky130_fd_sc_hd__a2bb2o_4
X_25459_ _25461_/CLK _12117_/X HRESETn VGND VGND VPWR VPWR _12116_/A sky130_fd_sc_hd__dfrtp_4
X_18000_ _18000_/A _18000_/B _18000_/C VGND VGND VPWR VPWR _18006_/B sky130_fd_sc_hd__and3_4
X_15212_ _15212_/A _15211_/X VGND VGND VPWR VPWR _15212_/X sky130_fd_sc_hd__or2_4
X_12424_ _25443_/Q _12424_/B VGND VGND VPWR VPWR _12425_/C sky130_fd_sc_hd__or2_4
XFILLER_107_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25109__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16192_ _16192_/A VGND VGND VPWR VPWR _16217_/A sky130_fd_sc_hd__buf_2
XFILLER_138_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15143_ _15336_/C _24589_/Q _24973_/Q _15086_/Y VGND VGND VPWR VPWR _15143_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17993__A _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12355_ _13029_/A _24830_/Q _13029_/A _24830_/Q VGND VGND VPWR VPWR _12355_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12286_ _12199_/Y _12286_/B _12286_/C _12188_/A VGND VGND VPWR VPWR _12432_/A sky130_fd_sc_hd__or4_4
X_15074_ _15073_/Y _24578_/Q _15073_/Y _24578_/Q VGND VGND VPWR VPWR _15074_/X sky130_fd_sc_hd__a2bb2o_4
X_19951_ _19951_/A VGND VGND VPWR VPWR _19964_/A sky130_fd_sc_hd__inv_2
XFILLER_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22588__B1 _24853_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14025_ _14012_/A _14022_/Y _14025_/C _14025_/D VGND VGND VPWR VPWR _14026_/A sky130_fd_sc_hd__or4_4
X_18902_ _18901_/Y VGND VGND VPWR VPWR _18902_/X sky130_fd_sc_hd__buf_2
XANTENNA__19453__B1 _19407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19882_ _23574_/Q VGND VGND VPWR VPWR _19882_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16267__B1 _16266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18833_ _18833_/A _18830_/X _18831_/X _18833_/D VGND VGND VPWR VPWR _18833_/X sky130_fd_sc_hd__or4_4
XFILLER_122_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24744__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18764_ _18763_/X VGND VGND VPWR VPWR _24129_/D sky130_fd_sc_hd__inv_2
XFILLER_110_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15976_ _12190_/Y _15975_/X _15897_/X _15975_/X VGND VGND VPWR VPWR _15976_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17715_ _21192_/A VGND VGND VPWR VPWR _21663_/A sky130_fd_sc_hd__buf_2
XFILLER_76_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14927_ _14927_/A VGND VGND VPWR VPWR _14927_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18695_ _18672_/Y _18694_/X VGND VGND VPWR VPWR _18695_/X sky130_fd_sc_hd__or2_4
XFILLER_97_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17646_ _17642_/A _17639_/X _17646_/C VGND VGND VPWR VPWR _17646_/X sky130_fd_sc_hd__and3_4
XFILLER_64_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14858_ _14799_/C _14813_/X _14799_/C _14813_/X VGND VGND VPWR VPWR _14858_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12577__A2_N _24857_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13809_ _11865_/X VGND VGND VPWR VPWR _16720_/A sky130_fd_sc_hd__buf_2
XFILLER_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17577_ _17577_/A VGND VGND VPWR VPWR _17577_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14789_ _14659_/B VGND VGND VPWR VPWR _14789_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19316_ _19315_/Y _19312_/X _19291_/X _19312_/X VGND VGND VPWR VPWR _23771_/D sky130_fd_sc_hd__a2bb2o_4
X_16528_ _16528_/A VGND VGND VPWR VPWR _16528_/X sky130_fd_sc_hd__buf_2
XFILLER_31_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19247_ _19246_/Y _19244_/X _16867_/X _19244_/X VGND VGND VPWR VPWR _23795_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25532__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16459_ _16728_/A _16459_/B VGND VGND VPWR VPWR _16466_/A sky130_fd_sc_hd__nor2_4
X_19178_ _19178_/A VGND VGND VPWR VPWR _19178_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18129_ _18097_/A _18129_/B _18128_/X VGND VGND VPWR VPWR _18129_/X sky130_fd_sc_hd__and3_4
XANTENNA__22291__A2 _22288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_104_0_HCLK clkbuf_7_52_0_HCLK/X VGND VGND VPWR VPWR _24355_/CLK sky130_fd_sc_hd__clkbuf_1
X_21140_ _20530_/B VGND VGND VPWR VPWR _21140_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17732__A1_N _21491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_167_0_HCLK clkbuf_7_83_0_HCLK/X VGND VGND VPWR VPWR _23388_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_132_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21071_ _21071_/A VGND VGND VPWR VPWR _22464_/A sky130_fd_sc_hd__buf_2
XANTENNA__12840__A _25383_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20022_ _17708_/A _18287_/A _17730_/X _19971_/X VGND VGND VPWR VPWR _20023_/A sky130_fd_sc_hd__or4_4
XFILLER_113_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24485__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24830_ _24830_/CLK _24830_/D HRESETn VGND VGND VPWR VPWR _24830_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24414__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24761_ _24830_/CLK _15947_/X HRESETn VGND VGND VPWR VPWR _24761_/Q sky130_fd_sc_hd__dfrtp_4
X_21973_ _24187_/Q _21985_/B VGND VGND VPWR VPWR _21973_/X sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_2_0_0_HCLK_A clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13492__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22751__B1 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23712_ _24930_/CLK _19481_/X VGND VGND VPWR VPWR _19480_/A sky130_fd_sc_hd__dfxtp_4
X_20924_ _20909_/X _20923_/Y _24490_/Q _20913_/X VGND VGND VPWR VPWR _24053_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24692_ _24692_/CLK _24692_/D HRESETn VGND VGND VPWR VPWR _16105_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_70_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16430__B1 _16143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _20855_/A VGND VGND VPWR VPWR _24037_/D sky130_fd_sc_hd__inv_2
XFILLER_54_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23643_ _23649_/CLK _19688_/X VGND VGND VPWR VPWR _13237_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22503__B1 _21587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20786_ _13136_/A VGND VGND VPWR VPWR _20786_/Y sky130_fd_sc_hd__inv_2
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23574_ _23550_/CLK _19883_/X VGND VGND VPWR VPWR _23574_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25313_ _23904_/CLK _13464_/X HRESETn VGND VGND VPWR VPWR _25313_/Q sky130_fd_sc_hd__dfrtp_4
X_22525_ _22421_/X VGND VGND VPWR VPWR _22525_/X sky130_fd_sc_hd__buf_2
XANTENNA__25273__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25202__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25244_ _25070_/CLK _25244_/D HRESETn VGND VGND VPWR VPWR _13565_/A sky130_fd_sc_hd__dfrtp_4
X_22456_ _21408_/A VGND VGND VPWR VPWR _23126_/A sky130_fd_sc_hd__buf_2
XFILLER_10_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_63_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21407_ _21320_/X _21407_/B _21361_/X _21407_/D VGND VGND VPWR VPWR _21407_/X sky130_fd_sc_hd__or4_4
X_22387_ _22384_/Y _22385_/X _22386_/X _13557_/A _22506_/B VGND VGND VPWR VPWR _22387_/X
+ sky130_fd_sc_hd__a32o_4
X_25175_ _25172_/CLK _14269_/X HRESETn VGND VGND VPWR VPWR _14268_/A sky130_fd_sc_hd__dfrtp_4
X_12140_ _25461_/Q _12139_/Y _25461_/Q _12139_/Y VGND VGND VPWR VPWR _12140_/X sky130_fd_sc_hd__a2bb2o_4
X_21338_ _14220_/A VGND VGND VPWR VPWR _21338_/X sky130_fd_sc_hd__buf_2
XANTENNA__21490__B1 _18299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24126_ _24133_/CLK _18777_/X HRESETn VGND VGND VPWR VPWR _24126_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12071_ _12071_/A VGND VGND VPWR VPWR _12072_/D sky130_fd_sc_hd__buf_2
X_21269_ _13593_/X VGND VGND VPWR VPWR _22505_/A sky130_fd_sc_hd__buf_2
XFILLER_85_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24057_ _24492_/CLK _20941_/X HRESETn VGND VGND VPWR VPWR _24057_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23008_ _23008_/A _21048_/B VGND VGND VPWR VPWR _23008_/X sky130_fd_sc_hd__or2_4
XFILLER_137_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15830_ _12318_/Y _15826_/X _15758_/X _15829_/X VGND VGND VPWR VPWR _24815_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20679__A _20678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15761_ _12542_/Y _15759_/X _15620_/X _15759_/X VGND VGND VPWR VPWR _24849_/D sky130_fd_sc_hd__a2bb2o_4
X_12973_ _12845_/A _12975_/B _12972_/Y VGND VGND VPWR VPWR _25358_/D sky130_fd_sc_hd__o21a_4
XANTENNA__13483__B1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24959_ _24957_/CLK _24959_/D HRESETn VGND VGND VPWR VPWR _13926_/C sky130_fd_sc_hd__dfrtp_4
X_17500_ _25517_/Q _17499_/Y _11759_/Y _24304_/Q VGND VGND VPWR VPWR _17505_/B sky130_fd_sc_hd__a2bb2o_4
X_14712_ _14712_/A VGND VGND VPWR VPWR _14712_/X sky130_fd_sc_hd__buf_2
X_11924_ _11924_/A _11899_/Y VGND VGND VPWR VPWR _11924_/X sky130_fd_sc_hd__and2_4
X_18480_ _18457_/Y _18479_/X VGND VGND VPWR VPWR _18490_/B sky130_fd_sc_hd__or2_4
X_15692_ _15677_/A _15685_/A VGND VGND VPWR VPWR _18019_/A sky130_fd_sc_hd__or2_4
XFILLER_72_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18410__B2 _18460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17431_ _24315_/Q VGND VGND VPWR VPWR _17431_/Y sky130_fd_sc_hd__inv_2
X_14643_ _14638_/X VGND VGND VPWR VPWR _14643_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17988__A _17996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11855_ _25509_/Q VGND VGND VPWR VPWR _11855_/Y sky130_fd_sc_hd__inv_2
X_17362_ _17370_/A _17360_/X _17362_/C VGND VGND VPWR VPWR _24337_/D sky130_fd_sc_hd__and3_4
X_14574_ _14558_/X _14579_/B _13568_/X _25084_/Q VGND VGND VPWR VPWR _14574_/X sky130_fd_sc_hd__and4_4
X_11786_ _11783_/Y _11777_/X _11784_/X _11785_/X VGND VGND VPWR VPWR _11786_/X sky130_fd_sc_hd__a2bb2o_4
X_19101_ _21382_/B _19098_/X _16888_/X _19098_/X VGND VGND VPWR VPWR _19101_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11797__B1 _11796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16313_ _22940_/A VGND VGND VPWR VPWR _16313_/Y sky130_fd_sc_hd__inv_2
X_13525_ _25293_/Q _20955_/B _13524_/X VGND VGND VPWR VPWR _25293_/D sky130_fd_sc_hd__a21o_4
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17293_ _17293_/A _17293_/B VGND VGND VPWR VPWR _17293_/X sky130_fd_sc_hd__or2_4
X_19032_ _19032_/A VGND VGND VPWR VPWR _19032_/Y sky130_fd_sc_hd__inv_2
X_16244_ _22539_/A VGND VGND VPWR VPWR _16244_/Y sky130_fd_sc_hd__inv_2
X_13456_ _13317_/A _19747_/A VGND VGND VPWR VPWR _13457_/C sky130_fd_sc_hd__or2_4
XFILLER_103_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25129__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12407_ _25447_/Q _12407_/B VGND VGND VPWR VPWR _12409_/B sky130_fd_sc_hd__or2_4
X_16175_ _16167_/X _16170_/X _16175_/C _16175_/D VGND VGND VPWR VPWR _16176_/A sky130_fd_sc_hd__or4_4
X_13387_ _13387_/A _13387_/B VGND VGND VPWR VPWR _13387_/X sky130_fd_sc_hd__or2_4
XANTENNA__19674__B1 _19599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24996__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15126_ _15126_/A VGND VGND VPWR VPWR _15126_/Y sky130_fd_sc_hd__inv_2
X_12338_ _25340_/Q _24825_/Q _13054_/A _12337_/Y VGND VGND VPWR VPWR _12339_/D sky130_fd_sc_hd__o22a_4
XFILLER_138_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24925__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15057_ _15057_/A VGND VGND VPWR VPWR _15057_/Y sky130_fd_sc_hd__inv_2
X_19934_ _22246_/B _19931_/X _19615_/X _19931_/X VGND VGND VPWR VPWR _19934_/X sky130_fd_sc_hd__a2bb2o_4
X_12269_ _25426_/Q VGND VGND VPWR VPWR _12269_/Y sky130_fd_sc_hd__inv_2
X_14008_ _14007_/X _13989_/X _13990_/X _14040_/D VGND VGND VPWR VPWR _14009_/B sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_5_17_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19865_ _19865_/A VGND VGND VPWR VPWR _22328_/B sky130_fd_sc_hd__inv_2
XFILLER_96_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18816_ _18682_/A _18818_/B _18815_/Y VGND VGND VPWR VPWR _18816_/X sky130_fd_sc_hd__o21a_4
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19796_ _19796_/A VGND VGND VPWR VPWR _21375_/B sky130_fd_sc_hd__inv_2
XFILLER_83_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15959_ HWDATA[19] VGND VGND VPWR VPWR _15959_/X sky130_fd_sc_hd__buf_2
X_18747_ _18747_/A VGND VGND VPWR VPWR _18747_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18678_ _24117_/Q VGND VGND VPWR VPWR _18678_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17629_ _24299_/Q _17628_/Y VGND VGND VPWR VPWR _17629_/X sky130_fd_sc_hd__or2_4
X_20640_ _14238_/Y _20628_/X _20619_/X _20639_/X VGND VGND VPWR VPWR _20641_/A sky130_fd_sc_hd__a211o_4
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21213__A _21069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20571_ _20571_/A _20570_/Y _20571_/C VGND VGND VPWR VPWR _20571_/X sky130_fd_sc_hd__and3_4
XANTENNA__17912__B1 _14620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22310_ _17349_/A _22419_/A _25427_/Q _21062_/Y VGND VGND VPWR VPWR _22311_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23290_ _23128_/A _23289_/X VGND VGND VPWR VPWR _23299_/B sky130_fd_sc_hd__nor2_4
XFILLER_34_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22241_ _21469_/A _22233_/X _22240_/X VGND VGND VPWR VPWR _22241_/X sky130_fd_sc_hd__and3_4
XFILLER_121_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18522__A _16448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22172_ _22172_/A _22172_/B VGND VGND VPWR VPWR _22172_/X sky130_fd_sc_hd__and2_4
XANTENNA__22044__A _21504_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24666__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21123_ _14430_/Y _14220_/A _21121_/Y _21335_/A VGND VGND VPWR VPWR _21123_/X sky130_fd_sc_hd__o22a_4
XFILLER_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16042__A _16042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21054_ _24701_/Q _15654_/A _21031_/X _21053_/X VGND VGND VPWR VPWR _21054_/X sky130_fd_sc_hd__a211o_4
XFILLER_99_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20005_ _22243_/B _20002_/X _19978_/X _20002_/X VGND VGND VPWR VPWR _23531_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22698__B _22298_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19353__A _17945_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_5_0_HCLK clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24813_ _24813_/CLK _24813_/D HRESETn VGND VGND VPWR VPWR _12296_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21527__A1 _16640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12268__B2 _24739_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21527__B2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24744_ _24792_/CLK _24744_/D HRESETn VGND VGND VPWR VPWR _22465_/A sky130_fd_sc_hd__dfrtp_4
X_21956_ _18230_/A _21955_/X VGND VGND VPWR VPWR _21956_/Y sky130_fd_sc_hd__nand2_4
XFILLER_70_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _24049_/Q _20901_/A _20906_/X VGND VGND VPWR VPWR _20907_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24675_ _24346_/CLK _24675_/D HRESETn VGND VGND VPWR VPWR _22395_/A sky130_fd_sc_hd__dfrtp_4
X_21887_ _21249_/A VGND VGND VPWR VPWR _21887_/X sky130_fd_sc_hd__buf_2
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17601__A _17885_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14965__B1 _25005_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ _23598_/CLK _23626_/D VGND VGND VPWR VPWR _13288_/B sky130_fd_sc_hd__dfxtp_4
X_20838_ _20837_/Y _20832_/Y _13658_/B VGND VGND VPWR VPWR _20838_/X sky130_fd_sc_hd__o21a_4
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11779__B1 _11778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16250__A1_N _16249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23557_ _25055_/CLK _23557_/D VGND VGND VPWR VPWR _23557_/Q sky130_fd_sc_hd__dfxtp_4
X_20769_ _20743_/X _20768_/Y _15587_/A _20747_/X VGND VGND VPWR VPWR _20769_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _13310_/A _13310_/B VGND VGND VPWR VPWR _13313_/B sky130_fd_sc_hd__or2_4
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22508_ _22505_/X _22506_/X _21950_/A _22507_/Y VGND VGND VPWR VPWR _22508_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14290_ _13527_/B _12026_/X _13524_/B VGND VGND VPWR VPWR _14291_/D sky130_fd_sc_hd__or3_4
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23488_ _23453_/CLK _20116_/X VGND VGND VPWR VPWR _20115_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13241_ _13248_/A VGND VGND VPWR VPWR _13320_/A sky130_fd_sc_hd__buf_2
X_25227_ _23967_/CLK _14068_/X HRESETn VGND VGND VPWR VPWR _25227_/Q sky130_fd_sc_hd__dfrtp_4
X_22439_ _21306_/X VGND VGND VPWR VPWR _22440_/C sky130_fd_sc_hd__buf_2
XANTENNA__19528__A _19528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19656__B1 _19462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13172_ _13191_/A _13172_/B _13171_/X VGND VGND VPWR VPWR _13172_/X sky130_fd_sc_hd__and3_4
X_25158_ _25305_/CLK _25158_/D HRESETn VGND VGND VPWR VPWR _25158_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12123_ _25456_/Q VGND VGND VPWR VPWR _12123_/Y sky130_fd_sc_hd__inv_2
X_24109_ _24109_/CLK _24109_/D HRESETn VGND VGND VPWR VPWR _20974_/B sky130_fd_sc_hd__dfstp_4
X_17980_ _17980_/A VGND VGND VPWR VPWR _18224_/A sky130_fd_sc_hd__buf_2
XFILLER_97_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24336__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_150_0_HCLK clkbuf_7_75_0_HCLK/X VGND VGND VPWR VPWR _24248_/CLK sky130_fd_sc_hd__clkbuf_1
X_25089_ _25093_/CLK _14533_/X HRESETn VGND VGND VPWR VPWR _21119_/A sky130_fd_sc_hd__dfrtp_4
X_12054_ _12054_/A VGND VGND VPWR VPWR _12054_/X sky130_fd_sc_hd__buf_2
X_16931_ _16130_/Y _24259_/Q _16130_/Y _24259_/Q VGND VGND VPWR VPWR _16932_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16862_ _19780_/A VGND VGND VPWR VPWR _16862_/Y sky130_fd_sc_hd__inv_2
X_19650_ _13356_/B VGND VGND VPWR VPWR _19650_/Y sky130_fd_sc_hd__inv_2
X_15813_ _12315_/Y _15809_/X _11784_/X _15812_/X VGND VGND VPWR VPWR _24826_/D sky130_fd_sc_hd__a2bb2o_4
X_18601_ _18601_/A VGND VGND VPWR VPWR _18782_/A sky130_fd_sc_hd__inv_2
X_19581_ _13787_/A _19581_/B _13777_/A _15662_/D VGND VGND VPWR VPWR _21143_/A sky130_fd_sc_hd__or4_4
X_16793_ _16792_/Y _16730_/A _16720_/X _16730_/A VGND VGND VPWR VPWR _16793_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22715__B1 _24821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18532_ _18464_/C _18532_/B VGND VGND VPWR VPWR _18542_/B sky130_fd_sc_hd__or2_4
XFILLER_133_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15744_ _15728_/X _15742_/X _15743_/X _24857_/Q _15740_/X VGND VGND VPWR VPWR _15744_/X
+ sky130_fd_sc_hd__a32o_4
X_12956_ _12964_/A _12956_/B _12956_/C VGND VGND VPWR VPWR _25364_/D sky130_fd_sc_hd__and3_4
XANTENNA__21017__B _21017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17198__B2 _17350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23971__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11907_ _11872_/X _11905_/X _11896_/X _11904_/Y VGND VGND VPWR VPWR _11907_/X sky130_fd_sc_hd__a2bb2o_4
X_18463_ _24159_/Q VGND VGND VPWR VPWR _18464_/D sky130_fd_sc_hd__inv_2
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25195__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15675_ _16640_/B _15674_/X VGND VGND VPWR VPWR _15675_/X sky130_fd_sc_hd__or2_4
X_12887_ _12887_/A _12886_/X VGND VGND VPWR VPWR _12887_/X sky130_fd_sc_hd__or2_4
XANTENNA__15748__A2 _15742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17414_ _21355_/A VGND VGND VPWR VPWR _17415_/A sky130_fd_sc_hd__buf_2
X_14626_ _14626_/A VGND VGND VPWR VPWR _21962_/A sky130_fd_sc_hd__inv_2
XFILLER_60_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11838_ _11838_/A VGND VGND VPWR VPWR _11838_/X sky130_fd_sc_hd__buf_2
X_18394_ _22154_/A _18393_/Y _16197_/Y _24172_/Q VGND VGND VPWR VPWR _18394_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22129__A _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17345_ _17246_/B VGND VGND VPWR VPWR _17350_/B sky130_fd_sc_hd__buf_2
X_14557_ _14586_/A VGND VGND VPWR VPWR _14557_/X sky130_fd_sc_hd__buf_2
X_11769_ _11766_/Y _11760_/X _11767_/X _11768_/X VGND VGND VPWR VPWR _25531_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22494__A2 _22442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15031__A _25005_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13508_ _12000_/Y _13507_/X _11847_/X _13507_/X VGND VGND VPWR VPWR _25298_/D sky130_fd_sc_hd__a2bb2o_4
X_17276_ _23246_/A _17276_/B VGND VGND VPWR VPWR _17278_/B sky130_fd_sc_hd__or2_4
X_14488_ _14481_/A VGND VGND VPWR VPWR _14488_/X sky130_fd_sc_hd__buf_2
X_19015_ _19014_/X VGND VGND VPWR VPWR _19030_/A sky130_fd_sc_hd__inv_2
XFILLER_31_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16227_ _22733_/A VGND VGND VPWR VPWR _16227_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13439_ _13173_/X _13435_/X _13438_/X VGND VGND VPWR VPWR _13439_/X sky130_fd_sc_hd__or3_4
XANTENNA__15966__A _15795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12195__B1 _25447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16158_ _16156_/Y _16152_/X _15471_/X _16157_/X VGND VGND VPWR VPWR _24672_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15109_ _24596_/Q VGND VGND VPWR VPWR _15109_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16089_ _16083_/Y _16088_/X _11743_/X _16088_/X VGND VGND VPWR VPWR _16089_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12390__A _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24077__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19917_ _22076_/B _19911_/X _19783_/X _19916_/X VGND VGND VPWR VPWR _23562_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24006__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22954__B1 _12366_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18622__A1 _24526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19848_ _19843_/Y _19847_/X _19777_/X _19847_/X VGND VGND VPWR VPWR _23588_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19779_ _23611_/Q VGND VGND VPWR VPWR _22215_/B sky130_fd_sc_hd__inv_2
XFILLER_7_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21509__A1 _21494_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21810_ _21650_/A _21810_/B VGND VGND VPWR VPWR _21812_/B sky130_fd_sc_hd__or2_4
XFILLER_3_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22790_ _22790_/A VGND VGND VPWR VPWR _22790_/X sky130_fd_sc_hd__buf_2
XFILLER_64_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21741_ _21741_/A _21741_/B VGND VGND VPWR VPWR _21741_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17421__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24460_ _25010_/CLK _16738_/X HRESETn VGND VGND VPWR VPWR _15015_/A sky130_fd_sc_hd__dfrtp_4
X_21672_ _21666_/X _21671_/X _21481_/X VGND VGND VPWR VPWR _21672_/X sky130_fd_sc_hd__o21a_4
XFILLER_52_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_26_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23411_ _24209_/CLK _23411_/D VGND VGND VPWR VPWR _22389_/A sky130_fd_sc_hd__dfxtp_4
X_20623_ _20623_/A VGND VGND VPWR VPWR _23972_/D sky130_fd_sc_hd__inv_2
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24391_ _24391_/CLK _17054_/X HRESETn VGND VGND VPWR VPWR _24391_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20554_ _14439_/Y _20533_/X _20547_/X _20553_/X VGND VGND VPWR VPWR _20554_/X sky130_fd_sc_hd__a211o_4
XFILLER_138_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23342_ _23342_/A _23341_/X VGND VGND VPWR VPWR _23342_/X sky130_fd_sc_hd__and2_4
XANTENNA__22890__C1 _22889_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24847__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14175__A1 _14169_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20485_ _14278_/A _20485_/B _20488_/B VGND VGND VPWR VPWR _20491_/A sky130_fd_sc_hd__and3_4
X_23273_ _21863_/X _23272_/X _22466_/X _24872_/Q _23102_/X VGND VGND VPWR VPWR _23274_/B
+ sky130_fd_sc_hd__a32o_4
X_25012_ _25016_/CLK _25012_/D HRESETn VGND VGND VPWR VPWR _15227_/A sky130_fd_sc_hd__dfrtp_4
X_22224_ _21260_/X _22204_/X _22219_/X _22222_/Y _22223_/X VGND VGND VPWR VPWR _22224_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_106_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22155_ _24540_/Q _21293_/X _21326_/X VGND VGND VPWR VPWR _22155_/X sky130_fd_sc_hd__o21a_4
X_21106_ _22988_/A VGND VGND VPWR VPWR _21106_/X sky130_fd_sc_hd__buf_2
XFILLER_120_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_223_0_HCLK clkbuf_8_223_0_HCLK/A VGND VGND VPWR VPWR _25010_/CLK sky130_fd_sc_hd__clkbuf_1
X_22086_ _14945_/A _21858_/X _21556_/X _22085_/X VGND VGND VPWR VPWR _22086_/X sky130_fd_sc_hd__a211o_4
XFILLER_134_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21037_ _21112_/B VGND VGND VPWR VPWR _21038_/B sky130_fd_sc_hd__inv_2
XFILLER_86_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23317__B _16795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16624__B1 _14555_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21118__A _21143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12810_ _12810_/A VGND VGND VPWR VPWR _12850_/B sky130_fd_sc_hd__inv_2
X_13790_ _14406_/A _21027_/B VGND VGND VPWR VPWR _14255_/A sky130_fd_sc_hd__or2_4
XANTENNA__12110__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22988_ _22988_/A VGND VGND VPWR VPWR _22988_/X sky130_fd_sc_hd__buf_2
XFILLER_43_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12459__B _13008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12741_ _21005_/A _12394_/X _12740_/Y VGND VGND VPWR VPWR _25387_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_1_0_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_0_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24727_ _24712_/CLK _24727_/D HRESETn VGND VGND VPWR VPWR _24727_/Q sky130_fd_sc_hd__dfrtp_4
X_21939_ _21454_/A _21937_/X _21938_/X VGND VGND VPWR VPWR _21939_/X sky130_fd_sc_hd__and3_4
X_15460_ _14280_/X _24069_/Q _15441_/Y _13893_/B _15434_/X VGND VGND VPWR VPWR _15460_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_70_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12672_ _12611_/B _12666_/X _12648_/A _12669_/B VGND VGND VPWR VPWR _12672_/X sky130_fd_sc_hd__a211o_4
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24658_ _24654_/CLK _24658_/D HRESETn VGND VGND VPWR VPWR _23068_/A sky130_fd_sc_hd__dfrtp_4
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _16057_/A VGND VGND VPWR VPWR _14411_/X sky130_fd_sc_hd__buf_2
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ _23609_/CLK _19788_/X VGND VGND VPWR VPWR _19786_/A sky130_fd_sc_hd__dfxtp_4
X_15391_ _15406_/A _15390_/X VGND VGND VPWR VPWR _15408_/A sky130_fd_sc_hd__or2_4
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12475__A _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24589_ _24984_/CLK _16399_/X HRESETn VGND VGND VPWR VPWR _24589_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ _17130_/A _17130_/B VGND VGND VPWR VPWR _17151_/A sky130_fd_sc_hd__or2_4
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _25152_/Q _14341_/Y _24094_/Q VGND VGND VPWR VPWR _14342_/X sky130_fd_sc_hd__o21a_4
XFILLER_7_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24588__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17061_ _17061_/A VGND VGND VPWR VPWR _17061_/Y sky130_fd_sc_hd__inv_2
X_14273_ _14273_/A VGND VGND VPWR VPWR _14273_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15363__B1 _15339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24517__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16012_ _16012_/A VGND VGND VPWR VPWR _16012_/Y sky130_fd_sc_hd__inv_2
X_13224_ _13233_/A VGND VGND VPWR VPWR _13450_/A sky130_fd_sc_hd__buf_2
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_33_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_67_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_3_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13155_ _24191_/Q VGND VGND VPWR VPWR _13155_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12106_ _25463_/Q VGND VGND VPWR VPWR _12106_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13086_ _13092_/A _13092_/B VGND VGND VPWR VPWR _13086_/X sky130_fd_sc_hd__or2_4
X_17963_ _17960_/X VGND VGND VPWR VPWR _17963_/X sky130_fd_sc_hd__buf_2
XFILLER_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19702_ _19702_/A VGND VGND VPWR VPWR _19702_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12037_ _12036_/Y _12034_/X _25478_/Q _12034_/X VGND VGND VPWR VPWR _25479_/D sky130_fd_sc_hd__a2bb2o_4
X_16914_ _24264_/Q VGND VGND VPWR VPWR _16914_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17894_ _17893_/Y _17889_/X _17893_/A _17891_/Y VGND VGND VPWR VPWR _17894_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16410__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16615__B1 _16355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19633_ _19631_/Y _19628_/X _19632_/X _19628_/X VGND VGND VPWR VPWR _19633_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21028__A _21028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25376__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16845_ _14890_/Y _16844_/X _16525_/X _16844_/X VGND VGND VPWR VPWR _16845_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19721__A _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25305__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16776_ _24440_/Q VGND VGND VPWR VPWR _16776_/Y sky130_fd_sc_hd__inv_2
X_19564_ _23683_/Q VGND VGND VPWR VPWR _22229_/B sky130_fd_sc_hd__inv_2
X_13988_ _14003_/A VGND VGND VPWR VPWR _14023_/A sky130_fd_sc_hd__buf_2
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15727_ _12539_/Y _15721_/X _11767_/X _15721_/X VGND VGND VPWR VPWR _15727_/X sky130_fd_sc_hd__a2bb2o_4
X_18515_ _18508_/X VGND VGND VPWR VPWR _18519_/B sky130_fd_sc_hd__inv_2
XANTENNA__23243__A _24563_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12939_ _12979_/A VGND VGND VPWR VPWR _12964_/A sky130_fd_sc_hd__buf_2
X_19495_ _19494_/Y VGND VGND VPWR VPWR _19495_/X sky130_fd_sc_hd__buf_2
XFILLER_94_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21911__A1 _21895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15658_ _15658_/A VGND VGND VPWR VPWR _15777_/B sky130_fd_sc_hd__buf_2
X_18446_ _16189_/Y _18455_/A _16189_/Y _18455_/A VGND VGND VPWR VPWR _18446_/X sky130_fd_sc_hd__a2bb2o_4
X_14609_ _14561_/X _14608_/Y _14557_/X _14602_/X _13566_/A VGND VGND VPWR VPWR _25072_/D
+ sky130_fd_sc_hd__a32o_4
X_18377_ _18377_/A VGND VGND VPWR VPWR _18377_/X sky130_fd_sc_hd__buf_2
X_15589_ _15587_/Y _15588_/X _11781_/X _15588_/X VGND VGND VPWR VPWR _15589_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12385__A _12385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17328_ _17327_/X VGND VGND VPWR VPWR _24344_/D sky130_fd_sc_hd__inv_2
Xclkbuf_7_115_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_230_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17259_ _17178_/Y _17282_/B VGND VGND VPWR VPWR _17260_/B sky130_fd_sc_hd__or2_4
XANTENNA__24258__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20270_ _20270_/A VGND VGND VPWR VPWR _21252_/B sky130_fd_sc_hd__inv_2
XFILLER_118_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16854__B1 _16717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17416__A _17416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23960_ _24069_/CLK _23960_/D HRESETn VGND VGND VPWR VPWR _20488_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_116_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_53_0_HCLK clkbuf_8_53_0_HCLK/A VGND VGND VPWR VPWR _24368_/CLK sky130_fd_sc_hd__clkbuf_1
X_22911_ _21306_/X VGND VGND VPWR VPWR _23117_/C sky130_fd_sc_hd__buf_2
XFILLER_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23891_ _25488_/CLK _18970_/X VGND VGND VPWR VPWR _23891_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25046__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22842_ _22714_/X _22842_/B VGND VGND VPWR VPWR _22842_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22155__A1 _24540_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22695__C _22695_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20166__B1 _20123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22773_ _22772_/X VGND VGND VPWR VPWR _22773_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18247__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24512_ _24561_/CLK _16598_/X HRESETn VGND VGND VPWR VPWR _16597_/A sky130_fd_sc_hd__dfrtp_4
X_21724_ _13509_/Y _21561_/X _12038_/Y _21562_/X VGND VGND VPWR VPWR _21724_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25492_ _23533_/CLK _25492_/D HRESETn VGND VGND VPWR VPWR _19992_/A sky130_fd_sc_hd__dfrtp_4
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24443_ _25002_/CLK _16772_/X HRESETn VGND VGND VPWR VPWR _15023_/A sky130_fd_sc_hd__dfrtp_4
X_21655_ _21459_/A _20013_/Y VGND VGND VPWR VPWR _21656_/C sky130_fd_sc_hd__or2_4
XANTENNA__21115__C1 _21114_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20606_ _23969_/Q _17404_/A VGND VGND VPWR VPWR _20606_/X sky130_fd_sc_hd__and2_4
X_24374_ _24391_/CLK _17117_/Y HRESETn VGND VGND VPWR VPWR _24374_/Q sky130_fd_sc_hd__dfrtp_4
X_21586_ _21741_/A _21586_/B VGND VGND VPWR VPWR _21586_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24681__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23325_ _16541_/A _22467_/X _22834_/X _23324_/X VGND VGND VPWR VPWR _23326_/C sky130_fd_sc_hd__a211o_4
X_20537_ _20537_/A _20537_/B VGND VGND VPWR VPWR _20537_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24610__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20468_ _20468_/A VGND VGND VPWR VPWR _20468_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23256_ _24596_/Q _23082_/B VGND VGND VPWR VPWR _23256_/X sky130_fd_sc_hd__or2_4
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22207_ _22078_/X _22207_/B _22206_/X VGND VGND VPWR VPWR _22207_/X sky130_fd_sc_hd__and3_4
XANTENNA__22091__B1 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18834__A1 _24550_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20399_ _20399_/A VGND VGND VPWR VPWR _20399_/Y sky130_fd_sc_hd__inv_2
X_23187_ _23187_/A _23310_/B VGND VGND VPWR VPWR _23187_/X sky130_fd_sc_hd__or2_4
XANTENNA__18861__A1_N _16457_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16845__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22138_ _22138_/A VGND VGND VPWR VPWR _22466_/A sky130_fd_sc_hd__buf_2
XANTENNA__12270__A2_N _22267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14960_ _15233_/A VGND VGND VPWR VPWR _14960_/Y sky130_fd_sc_hd__inv_2
X_22069_ _21624_/A _22067_/X _22069_/C VGND VGND VPWR VPWR _22069_/X sky130_fd_sc_hd__and3_4
XFILLER_134_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18598__B1 _16594_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13911_ _13895_/X _13897_/X _13918_/A _13898_/Y VGND VGND VPWR VPWR _13911_/X sky130_fd_sc_hd__o22a_4
XFILLER_47_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14891_ _25022_/Q VGND VGND VPWR VPWR _15187_/A sky130_fd_sc_hd__inv_2
XFILLER_59_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16630_ _16630_/A VGND VGND VPWR VPWR _16630_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13842_ _13549_/Y _13839_/X _13797_/X _13839_/X VGND VGND VPWR VPWR _13842_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16561_ _16560_/Y _16558_/X _16300_/X _16558_/X VGND VGND VPWR VPWR _24527_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13773_ _24065_/Q VGND VGND VPWR VPWR _16725_/B sky130_fd_sc_hd__buf_2
XFILLER_90_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20157__B1 _20089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15512_ _15510_/Y _15511_/X HADDR[14] _15511_/X VGND VGND VPWR VPWR _24926_/D sky130_fd_sc_hd__a2bb2o_4
X_18300_ _18300_/A VGND VGND VPWR VPWR _18303_/B sky130_fd_sc_hd__inv_2
X_12724_ _12560_/A _12724_/B VGND VGND VPWR VPWR _12725_/B sky130_fd_sc_hd__or2_4
X_19280_ _23782_/Q VGND VGND VPWR VPWR _21381_/B sky130_fd_sc_hd__inv_2
XFILLER_91_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16492_ _16490_/Y _16486_/X _16405_/X _16491_/X VGND VGND VPWR VPWR _16492_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24769__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18231_ _18231_/A VGND VGND VPWR VPWR _18249_/A sky130_fd_sc_hd__inv_2
XFILLER_130_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15443_ _13919_/X _15437_/X _15432_/X _13956_/A _15438_/X VGND VGND VPWR VPWR _24958_/D
+ sky130_fd_sc_hd__a32o_4
X_12655_ _12517_/Y _12652_/X _12654_/Y VGND VGND VPWR VPWR _12655_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15584__B1 _11774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17996__A _17996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18162_ _15694_/X _18146_/X _18161_/X _24232_/Q _18019_/X VGND VGND VPWR VPWR _18162_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15374_ _15374_/A _15373_/Y VGND VGND VPWR VPWR _15375_/C sky130_fd_sc_hd__or2_4
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ _24864_/Q VGND VGND VPWR VPWR _12586_/Y sky130_fd_sc_hd__inv_2
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17113_ _17100_/X VGND VGND VPWR VPWR _17114_/B sky130_fd_sc_hd__inv_2
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ _14325_/A VGND VGND VPWR VPWR _14325_/X sky130_fd_sc_hd__buf_2
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18093_ _18054_/X _23817_/Q VGND VGND VPWR VPWR _18095_/B sky130_fd_sc_hd__or2_4
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24351__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16405__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17044_ _17130_/A _17044_/B _16993_/Y _17043_/Y VGND VGND VPWR VPWR _17045_/C sky130_fd_sc_hd__or4_4
X_14256_ _21139_/B VGND VGND VPWR VPWR _14257_/A sky130_fd_sc_hd__buf_2
X_13207_ _13413_/A _13204_/X _13206_/X VGND VGND VPWR VPWR _13207_/X sky130_fd_sc_hd__and3_4
X_14187_ _12052_/B VGND VGND VPWR VPWR _15549_/B sky130_fd_sc_hd__inv_2
XFILLER_87_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22621__A2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18829__A1_N _16476_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15639__B2 _15563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13138_ _24028_/Q _13137_/X VGND VGND VPWR VPWR _20675_/B sky130_fd_sc_hd__or2_4
X_18995_ _18995_/A VGND VGND VPWR VPWR _18995_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13069_ _13068_/X VGND VGND VPWR VPWR _13069_/Y sky130_fd_sc_hd__inv_2
X_17946_ _17930_/A _17946_/B VGND VGND VPWR VPWR _17947_/C sky130_fd_sc_hd__or2_4
XFILLER_26_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16140__A _22556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17877_ _16927_/X _17848_/B VGND VGND VPWR VPWR _17878_/B sky130_fd_sc_hd__or2_4
XFILLER_26_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19616_ _19614_/Y _19611_/X _19615_/X _19611_/X VGND VGND VPWR VPWR _23667_/D sky130_fd_sc_hd__a2bb2o_4
X_16828_ _16827_/Y _16825_/X _15743_/X _16825_/X VGND VGND VPWR VPWR _16828_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19547_ _15766_/A VGND VGND VPWR VPWR _19547_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16759_ _16773_/A VGND VGND VPWR VPWR _16759_/X sky130_fd_sc_hd__buf_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19478_ _23713_/Q VGND VGND VPWR VPWR _21941_/B sky130_fd_sc_hd__inv_2
XFILLER_34_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18429_ _16237_/Y _24157_/Q _16237_/Y _24157_/Q VGND VGND VPWR VPWR _18429_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11731__B _13777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24439__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21440_ _15784_/B VGND VGND VPWR VPWR _22429_/A sky130_fd_sc_hd__buf_2
XANTENNA__21859__C _21859_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21371_ _21371_/A _19838_/Y VGND VGND VPWR VPWR _21374_/B sky130_fd_sc_hd__or2_4
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24092__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12843__A _12843_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20322_ _20317_/X _19586_/D _13835_/A _22389_/A _20326_/A VGND VGND VPWR VPWR _23411_/D
+ sky130_fd_sc_hd__a32o_4
X_23110_ _24693_/Q _22864_/X VGND VGND VPWR VPWR _23110_/X sky130_fd_sc_hd__or2_4
XANTENNA__24021__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24090_ _25246_/CLK _24090_/D HRESETn VGND VGND VPWR VPWR _12015_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_66_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20253_ _20252_/X VGND VGND VPWR VPWR _20266_/A sky130_fd_sc_hd__inv_2
XANTENNA__23223__A1_N _12385_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23041_ _22770_/X _23039_/X _23040_/X _24726_/Q _22972_/X VGND VGND VPWR VPWR _23041_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_89_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12281__C _12280_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20184_ _23462_/Q VGND VGND VPWR VPWR _20184_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25298__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23022__C1 _23021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25227__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24992_ _24984_/CLK _24992_/D HRESETn VGND VGND VPWR VPWR _15322_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23943_ _25205_/CLK _23943_/D HRESETn VGND VGND VPWR VPWR _23943_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20387__B1 _19758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23874_ _25485_/CLK _23874_/D VGND VGND VPWR VPWR _23874_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23325__B1 _22834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16602__A1_N _16599_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22825_ _20892_/Y _22824_/X _20754_/C _22280_/A VGND VGND VPWR VPWR _22825_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17004__B1 _24713_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22756_ _22739_/Y _22744_/Y _22752_/Y _21437_/X _22755_/X VGND VGND VPWR VPWR _22756_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24862__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21707_ _21275_/X _21693_/X _21696_/X _21703_/X _21706_/X VGND VGND VPWR VPWR _21707_/X
+ sky130_fd_sc_hd__o41a_4
XANTENNA__15566__B1 _11749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25475_ _25461_/CLK _25475_/D HRESETn VGND VGND VPWR VPWR _25475_/Q sky130_fd_sc_hd__dfrtp_4
X_22687_ _22687_/A VGND VGND VPWR VPWR _22719_/A sky130_fd_sc_hd__inv_2
XANTENNA__18705__A _18705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16617__A1_N _16616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12440_ _12199_/Y _12286_/B _12440_/C _12432_/B VGND VGND VPWR VPWR _12440_/X sky130_fd_sc_hd__or4_4
XFILLER_40_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24426_ _24457_/CLK _16810_/X HRESETn VGND VGND VPWR VPWR _16809_/A sky130_fd_sc_hd__dfrtp_4
X_21638_ _21995_/A VGND VGND VPWR VPWR _22390_/B sky130_fd_sc_hd__buf_2
XFILLER_90_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22300__A1 _14922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12371_ _12371_/A _12365_/X _12371_/C _12371_/D VGND VGND VPWR VPWR _12381_/C sky130_fd_sc_hd__or4_4
X_24357_ _24318_/CLK _17278_/X HRESETn VGND VGND VPWR VPWR _23246_/A sky130_fd_sc_hd__dfrtp_4
X_21569_ _21547_/Y _21555_/X _21558_/X _21568_/Y VGND VGND VPWR VPWR _21569_/X sky130_fd_sc_hd__a211o_4
XFILLER_5_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14110_ _14129_/A VGND VGND VPWR VPWR _14110_/X sky130_fd_sc_hd__buf_2
X_23308_ _21512_/X _23307_/X _21514_/X _24734_/Q _21520_/X VGND VGND VPWR VPWR _23308_/X
+ sky130_fd_sc_hd__a32o_4
X_15090_ _15090_/A VGND VGND VPWR VPWR _15090_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20970__A scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24288_ _24288_/CLK _24288_/D HRESETn VGND VGND VPWR VPWR _24288_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14041_ _14041_/A VGND VGND VPWR VPWR _14041_/Y sky130_fd_sc_hd__inv_2
X_23239_ _23207_/A _23236_/X _23239_/C VGND VGND VPWR VPWR _23240_/D sky130_fd_sc_hd__and3_4
XANTENNA__22603__A2 _22425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16818__B1 HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17800_ _17799_/X VGND VGND VPWR VPWR _17800_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17056__A _17384_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15992_ _16371_/A _15992_/B VGND VGND VPWR VPWR _16276_/B sky130_fd_sc_hd__or2_4
X_18780_ _18742_/A VGND VGND VPWR VPWR _18799_/A sky130_fd_sc_hd__buf_2
X_14943_ _15227_/A _14941_/Y _14942_/Y _14945_/A VGND VGND VPWR VPWR _14943_/X sky130_fd_sc_hd__a2bb2o_4
X_17731_ _17730_/X _17724_/A _17729_/A _17724_/Y VGND VGND VPWR VPWR _17731_/X sky130_fd_sc_hd__o22a_4
XFILLER_121_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15811__A1_N _12366_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14874_ _14868_/Y _14810_/X _14811_/X _14873_/X VGND VGND VPWR VPWR _14874_/X sky130_fd_sc_hd__o22a_4
X_17662_ _17662_/A _17662_/B _17578_/C _17695_/A VGND VGND VPWR VPWR _17662_/X sky130_fd_sc_hd__or4_4
XANTENNA__22119__A1 _13784_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19401_ _19401_/A VGND VGND VPWR VPWR _19401_/X sky130_fd_sc_hd__buf_2
XFILLER_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20393__A3 _11867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13825_ _13822_/A VGND VGND VPWR VPWR _13825_/X sky130_fd_sc_hd__buf_2
X_16613_ _24506_/Q VGND VGND VPWR VPWR _16613_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21306__A _21306_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17593_ _17611_/A _17583_/X VGND VGND VPWR VPWR _17604_/A sky130_fd_sc_hd__or2_4
XANTENNA__12928__A _12936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11832__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16544_ _16550_/A VGND VGND VPWR VPWR _16545_/A sky130_fd_sc_hd__buf_2
X_19332_ _14663_/D _18987_/D _19399_/C VGND VGND VPWR VPWR _19332_/X sky130_fd_sc_hd__or3_4
X_13756_ _13736_/X _13748_/X _20077_/A VGND VGND VPWR VPWR _13756_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_16_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12707_ _12707_/A _12707_/B VGND VGND VPWR VPWR _12708_/B sky130_fd_sc_hd__or2_4
X_16475_ _16473_/Y _16474_/X _16297_/X _16474_/X VGND VGND VPWR VPWR _16475_/X sky130_fd_sc_hd__a2bb2o_4
X_19263_ _13748_/C _13757_/B _13746_/A VGND VGND VPWR VPWR _19845_/C sky130_fd_sc_hd__or3_4
X_13687_ _13718_/A _13686_/X VGND VGND VPWR VPWR _13688_/B sky130_fd_sc_hd__or2_4
XANTENNA__24532__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15426_ _13953_/A _13947_/A _13930_/D VGND VGND VPWR VPWR _15426_/X sky130_fd_sc_hd__or3_4
X_18214_ _18150_/A _18214_/B VGND VGND VPWR VPWR _18214_/X sky130_fd_sc_hd__or2_4
X_12638_ _12524_/Y _12620_/X _12645_/A _12629_/X VGND VGND VPWR VPWR _12638_/X sky130_fd_sc_hd__or4_4
X_19194_ _19193_/Y _19188_/X _19149_/X _19175_/Y VGND VGND VPWR VPWR _19194_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13032__A1 _12299_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22137__A _16352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18334__B _17449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15357_ _15372_/A _15357_/B _15357_/C VGND VGND VPWR VPWR _15357_/X sky130_fd_sc_hd__and3_4
X_18145_ _18177_/A _18141_/X _18145_/C VGND VGND VPWR VPWR _18146_/C sky130_fd_sc_hd__or3_4
XFILLER_8_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ _12569_/A _12564_/X _12566_/X _12568_/X VGND VGND VPWR VPWR _12569_/X sky130_fd_sc_hd__or4_4
XFILLER_89_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14308_ MSO_S2 _14307_/X _25164_/Q _14302_/X VGND VGND VPWR VPWR _14308_/Y sky130_fd_sc_hd__a22oi_4
X_18076_ _18181_/A _18073_/X _18076_/C VGND VGND VPWR VPWR _18077_/C sky130_fd_sc_hd__and3_4
XFILLER_32_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15288_ _15246_/A _15248_/B _15287_/X VGND VGND VPWR VPWR _15288_/X sky130_fd_sc_hd__and3_4
X_17027_ _17085_/A VGND VGND VPWR VPWR _17048_/A sky130_fd_sc_hd__inv_2
X_14239_ _11862_/A VGND VGND VPWR VPWR _14239_/X sky130_fd_sc_hd__buf_2
XANTENNA__14532__A1 _21119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25391__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25320__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18978_ _18972_/A VGND VGND VPWR VPWR _18978_/X sky130_fd_sc_hd__buf_2
XFILLER_67_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17929_ _17929_/A _23876_/Q VGND VGND VPWR VPWR _17931_/B sky130_fd_sc_hd__or2_4
XANTENNA__11726__B _11726_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20940_ _24057_/Q _13666_/X _20939_/X VGND VGND VPWR VPWR _20940_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_82_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20384__A3 _11838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20871_ _24041_/Q _13662_/B _20870_/Y VGND VGND VPWR VPWR _20871_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_26_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15796__B1 _24837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_127_0_HCLK clkbuf_7_63_0_HCLK/X VGND VGND VPWR VPWR _24980_/CLK sky130_fd_sc_hd__clkbuf_1
X_22610_ _24413_/Q _22523_/X _22524_/X _22609_/X VGND VGND VPWR VPWR _22611_/C sky130_fd_sc_hd__a211o_4
XANTENNA__21869__B1 _24811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23590_ _24089_/CLK _19839_/X VGND VGND VPWR VPWR _19838_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_4_6_0_HCLK_A clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22541_ _24544_/Q _22422_/X _22527_/X VGND VGND VPWR VPWR _22541_/X sky130_fd_sc_hd__o21a_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24273__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25260_ _25070_/CLK _25260_/D HRESETn VGND VGND VPWR VPWR _13802_/A sky130_fd_sc_hd__dfrtp_4
X_22472_ _24781_/Q _22472_/B VGND VGND VPWR VPWR _22472_/X sky130_fd_sc_hd__or2_4
XANTENNA__24202__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24211_ _24214_/CLK _24211_/D HRESETn VGND VGND VPWR VPWR _24211_/Q sky130_fd_sc_hd__dfrtp_4
X_21423_ _21422_/X VGND VGND VPWR VPWR _23314_/B sky130_fd_sc_hd__buf_2
XFILLER_120_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25191_ _25192_/CLK _14213_/X HRESETn VGND VGND VPWR VPWR _14212_/A sky130_fd_sc_hd__dfrtp_4
X_24142_ _24136_/CLK _24142_/D HRESETn VGND VGND VPWR VPWR _24142_/Q sky130_fd_sc_hd__dfrtp_4
X_21354_ _25232_/Q VGND VGND VPWR VPWR _21354_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25479__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20305_ _22028_/B _20299_/X _19981_/X _20304_/X VGND VGND VPWR VPWR _23417_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15720__B1 _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25408__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24073_ _24117_/CLK _24073_/D HRESETn VGND VGND VPWR VPWR _24073_/Q sky130_fd_sc_hd__dfrtp_4
X_21285_ _21285_/A VGND VGND VPWR VPWR _21290_/C sky130_fd_sc_hd__buf_2
X_23024_ _22714_/X _23024_/B VGND VGND VPWR VPWR _23024_/Y sky130_fd_sc_hd__nor2_4
X_20236_ _20235_/Y _20233_/X _19755_/X _20233_/X VGND VGND VPWR VPWR _23443_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20167_ _23468_/Q VGND VGND VPWR VPWR _22376_/B sky130_fd_sc_hd__inv_2
XANTENNA__25061__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17307__C _17346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20098_ _23494_/Q VGND VGND VPWR VPWR _20098_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23010__A2 _21021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24975_ _24977_/CLK _15386_/Y HRESETn VGND VGND VPWR VPWR _24975_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22510__A _22510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11940_ _11938_/Y _11935_/X _11939_/X _11935_/X VGND VGND VPWR VPWR _25494_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23926_ _24077_/CLK _20979_/Y HRESETn VGND VGND VPWR VPWR _23926_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_72_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_23_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21572__A2 _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18973__B1 _17424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_86_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_86_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11871_ _11871_/A VGND VGND VPWR VPWR _11871_/Y sky130_fd_sc_hd__inv_2
X_23857_ _23854_/CLK _19072_/X VGND VGND VPWR VPWR _23857_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13610_ _13610_/A VGND VGND VPWR VPWR _18088_/A sky130_fd_sc_hd__buf_2
XANTENNA__11652__A _21504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22808_ _16452_/A VGND VGND VPWR VPWR _22808_/X sky130_fd_sc_hd__buf_2
X_14590_ _13769_/Y VGND VGND VPWR VPWR _14590_/X sky130_fd_sc_hd__buf_2
X_23788_ _24398_/CLK _19267_/X VGND VGND VPWR VPWR _23788_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13541_ _13541_/A _13541_/B _13541_/C VGND VGND VPWR VPWR _13541_/X sky130_fd_sc_hd__and3_4
XANTENNA__23115__A1_N _12277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25527_ _25436_/CLK _11782_/X HRESETn VGND VGND VPWR VPWR _25527_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15539__B1 HADDR[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22739_ _22549_/A _22738_/X VGND VGND VPWR VPWR _22739_/Y sky130_fd_sc_hd__nand2_4
XFILLER_71_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16260_ _16258_/Y _16254_/X _15471_/X _16259_/X VGND VGND VPWR VPWR _16260_/X sky130_fd_sc_hd__a2bb2o_4
X_13472_ _11867_/A VGND VGND VPWR VPWR _13472_/X sky130_fd_sc_hd__buf_2
X_25458_ _24097_/CLK _25458_/D HRESETn VGND VGND VPWR VPWR _25458_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14211__B1 _13803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14682__B _14682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15211_ _15211_/A _15211_/B VGND VGND VPWR VPWR _15211_/X sky130_fd_sc_hd__or2_4
XANTENNA__21088__A1 _24632_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12423_ _12414_/X VGND VGND VPWR VPWR _12424_/B sky130_fd_sc_hd__inv_2
XFILLER_51_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24409_ _24998_/CLK _16842_/X HRESETn VGND VGND VPWR VPWR _24409_/Q sky130_fd_sc_hd__dfrtp_4
X_16191_ _23242_/A VGND VGND VPWR VPWR _16191_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12483__A _12220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25389_ _25411_/CLK _25389_/D HRESETn VGND VGND VPWR VPWR _25389_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12773__B1 _12841_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19150__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23996__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15142_ _24985_/Q VGND VGND VPWR VPWR _15336_/C sky130_fd_sc_hd__inv_2
XFILLER_126_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12354_ _25345_/Q VGND VGND VPWR VPWR _13029_/A sky130_fd_sc_hd__inv_2
XANTENNA__21796__A _21658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23925__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15073_ _24974_/Q VGND VGND VPWR VPWR _15073_/Y sky130_fd_sc_hd__inv_2
X_19950_ _20338_/A _20338_/B _19492_/X VGND VGND VPWR VPWR _19951_/A sky130_fd_sc_hd__or3_4
XANTENNA__25149__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12285_ _12248_/Y _12238_/A _12285_/C _12433_/A VGND VGND VPWR VPWR _12285_/X sky130_fd_sc_hd__or4_4
XANTENNA__18170__A _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14024_ _14002_/X _13992_/X VGND VGND VPWR VPWR _14025_/D sky130_fd_sc_hd__or2_4
X_18901_ _18900_/X VGND VGND VPWR VPWR _18901_/Y sky130_fd_sc_hd__inv_2
X_19881_ _21650_/B _19880_/X _19629_/X _19880_/X VGND VGND VPWR VPWR _19881_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18832_ _16483_/Y _18658_/A _16483_/Y _18658_/A VGND VGND VPWR VPWR _18833_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18763_ _18753_/C _18756_/B _18733_/X _18760_/Y VGND VGND VPWR VPWR _18763_/X sky130_fd_sc_hd__a211o_4
XFILLER_23_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15975_ _15937_/Y VGND VGND VPWR VPWR _15975_/X sky130_fd_sc_hd__buf_2
XANTENNA__22420__A _22419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17714_ _24199_/Q VGND VGND VPWR VPWR _21192_/A sky130_fd_sc_hd__buf_2
XANTENNA__16509__A1_N _16508_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14926_ _15067_/C VGND VGND VPWR VPWR _14926_/X sky130_fd_sc_hd__buf_2
X_18694_ _18673_/Y _18658_/Y _18676_/X _18693_/X VGND VGND VPWR VPWR _18694_/X sky130_fd_sc_hd__or4_4
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24784__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18964__B1 _18940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21036__A _22835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17645_ _17564_/Y _17645_/B VGND VGND VPWR VPWR _17646_/C sky130_fd_sc_hd__nand2_4
X_14857_ _14843_/X _14856_/Y _14814_/C _14843_/X VGND VGND VPWR VPWR _14857_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24713__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13808_ _25258_/Q VGND VGND VPWR VPWR _13808_/Y sky130_fd_sc_hd__inv_2
X_14788_ _18017_/A _14667_/X _18017_/A _14667_/X VGND VGND VPWR VPWR _14792_/C sky130_fd_sc_hd__a2bb2o_4
X_17576_ _17576_/A VGND VGND VPWR VPWR _17576_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14450__B1 _14239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19315_ _17974_/B VGND VGND VPWR VPWR _19315_/Y sky130_fd_sc_hd__inv_2
X_13739_ _21643_/A _13739_/B VGND VGND VPWR VPWR _13744_/B sky130_fd_sc_hd__or2_4
X_16527_ _24539_/Q VGND VGND VPWR VPWR _16527_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19246_ _19246_/A VGND VGND VPWR VPWR _19246_/Y sky130_fd_sc_hd__inv_2
X_16458_ _15931_/B VGND VGND VPWR VPWR _16728_/A sky130_fd_sc_hd__buf_2
XANTENNA__14202__B1 _13835_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15409_ _15409_/A VGND VGND VPWR VPWR _15409_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16389_ _16389_/A VGND VGND VPWR VPWR _16389_/X sky130_fd_sc_hd__buf_2
X_19177_ _19173_/Y _19176_/X _19155_/X _19176_/X VGND VGND VPWR VPWR _19177_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15950__B1 _15949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18128_ _18058_/A _18128_/B _18127_/X VGND VGND VPWR VPWR _18128_/X sky130_fd_sc_hd__or3_4
X_18059_ _18059_/A _18059_/B _18058_/X VGND VGND VPWR VPWR _18059_/X sky130_fd_sc_hd__and3_4
XANTENNA__25501__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21070_ _23019_/B VGND VGND VPWR VPWR _23069_/B sky130_fd_sc_hd__buf_2
XFILLER_28_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20021_ _23524_/Q VGND VGND VPWR VPWR _22329_/B sky130_fd_sc_hd__inv_2
XFILLER_99_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11737__A _21582_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14269__B1 _13800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22907__A1_N _12286_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17424__A _16528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24760_ _24830_/CLK _15948_/X HRESETn VGND VGND VPWR VPWR _24760_/Q sky130_fd_sc_hd__dfrtp_4
X_21972_ _18365_/A _20335_/Y _24187_/Q _21985_/B VGND VGND VPWR VPWR _21972_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23711_ _23711_/CLK _23711_/D VGND VGND VPWR VPWR _23711_/Q sky130_fd_sc_hd__dfxtp_4
X_20923_ _24053_/Q _20922_/B _20922_/Y VGND VGND VPWR VPWR _20923_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__15769__B1 _24845_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24691_ _24691_/CLK _24691_/D HRESETn VGND VGND VPWR VPWR _23043_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24454__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23642_ _23649_/CLK _19691_/X VGND VGND VPWR VPWR _19689_/A sky130_fd_sc_hd__dfxtp_4
X_20854_ _16699_/Y _20836_/X _20845_/X _20853_/Y VGND VGND VPWR VPWR _20855_/A sky130_fd_sc_hd__o22a_4
XFILLER_78_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22503__A1 _13813_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23573_ _24309_/CLK _19886_/X VGND VGND VPWR VPWR _19884_/A sky130_fd_sc_hd__dfxtp_4
X_20785_ _20770_/X _20784_/Y _15577_/A _20774_/X VGND VGND VPWR VPWR _20785_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19380__B1 _19313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25312_ _24383_/CLK _13473_/X HRESETn VGND VGND VPWR VPWR _23343_/A sky130_fd_sc_hd__dfrtp_4
X_22524_ _22524_/A VGND VGND VPWR VPWR _22524_/X sky130_fd_sc_hd__buf_2
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16194__B1 _15940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14744__A1 _21781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25243_ _25070_/CLK _13847_/X HRESETn VGND VGND VPWR VPWR _13846_/A sky130_fd_sc_hd__dfrtp_4
X_22455_ _21588_/X VGND VGND VPWR VPWR _22783_/A sky130_fd_sc_hd__buf_2
XANTENNA__15941__B1 _15940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21406_ _21405_/X VGND VGND VPWR VPWR _21407_/D sky130_fd_sc_hd__inv_2
XFILLER_109_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25174_ _24883_/CLK _14272_/X HRESETn VGND VGND VPWR VPWR _25174_/Q sky130_fd_sc_hd__dfrtp_4
X_22386_ _22386_/A _22390_/B VGND VGND VPWR VPWR _22386_/X sky130_fd_sc_hd__or2_4
XANTENNA__22019__B1 _21679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24125_ _24133_/CLK _24125_/D HRESETn VGND VGND VPWR VPWR _18686_/A sky130_fd_sc_hd__dfrtp_4
X_21337_ _14177_/Y _22316_/B _23920_/Q _21351_/B VGND VGND VPWR VPWR _21343_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25242__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12070_ _16453_/B VGND VGND VPWR VPWR _12071_/A sky130_fd_sc_hd__buf_2
XFILLER_46_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24056_ _24055_/CLK _20937_/Y HRESETn VGND VGND VPWR VPWR _24056_/Q sky130_fd_sc_hd__dfrtp_4
X_21268_ _18270_/X _21266_/X _21162_/X _21267_/Y VGND VGND VPWR VPWR _21268_/X sky130_fd_sc_hd__a211o_4
XFILLER_1_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23007_ _22808_/X _23007_/B _23007_/C VGND VGND VPWR VPWR _23007_/X sky130_fd_sc_hd__and3_4
X_20219_ _23449_/Q VGND VGND VPWR VPWR _20219_/Y sky130_fd_sc_hd__inv_2
X_21199_ _19535_/X _21333_/A VGND VGND VPWR VPWR _21200_/B sky130_fd_sc_hd__or2_4
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23336__A _23336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19199__B1 _19155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15760_ _12536_/Y _15754_/X _15758_/X _15759_/X VGND VGND VPWR VPWR _15760_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12972_ _12845_/A _12975_/B _12866_/X VGND VGND VPWR VPWR _12972_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_131_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24958_ _24957_/CLK _24958_/D HRESETn VGND VGND VPWR VPWR _24958_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11923_ _19612_/A VGND VGND VPWR VPWR _11923_/Y sky130_fd_sc_hd__inv_2
X_14711_ _14710_/Y VGND VGND VPWR VPWR _14712_/A sky130_fd_sc_hd__buf_2
XFILLER_79_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15691_ _15690_/X VGND VGND VPWR VPWR _15691_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23909_ _23453_/CLK _23909_/D VGND VGND VPWR VPWR _23909_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24195__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24889_ _24889_/CLK _15615_/X HRESETn VGND VGND VPWR VPWR _15614_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_75_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14642_ _18059_/A _14641_/X _18059_/A _14641_/X VGND VGND VPWR VPWR _14642_/X sky130_fd_sc_hd__a2bb2o_4
X_17430_ _17429_/Y _17425_/X _16787_/X _17425_/X VGND VGND VPWR VPWR _24316_/D sky130_fd_sc_hd__a2bb2o_4
X_11854_ _11850_/Y _11848_/X _11853_/X _11848_/X VGND VGND VPWR VPWR _25510_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24124__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_110_0_HCLK clkbuf_7_55_0_HCLK/X VGND VGND VPWR VPWR _24889_/CLK sky130_fd_sc_hd__clkbuf_1
X_14573_ _14573_/A VGND VGND VPWR VPWR _14579_/B sky130_fd_sc_hd__inv_2
X_17361_ _17350_/A _17361_/B VGND VGND VPWR VPWR _17362_/C sky130_fd_sc_hd__or2_4
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15789__A _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11785_ _11777_/A VGND VGND VPWR VPWR _11785_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_173_0_HCLK clkbuf_7_86_0_HCLK/X VGND VGND VPWR VPWR _23533_/CLK sky130_fd_sc_hd__clkbuf_1
X_19100_ _19100_/A VGND VGND VPWR VPWR _21382_/B sky130_fd_sc_hd__inv_2
XANTENNA__19371__B1 _19370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13524_ _20953_/B _13524_/B VGND VGND VPWR VPWR _13524_/X sky130_fd_sc_hd__and2_4
X_16312_ _16310_/Y _16311_/X _15955_/X _16311_/X VGND VGND VPWR VPWR _24620_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17292_ _17257_/A _17291_/X VGND VGND VPWR VPWR _17293_/B sky130_fd_sc_hd__or2_4
XFILLER_14_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16243_ _16240_/Y _16241_/X _16242_/X _16241_/X VGND VGND VPWR VPWR _24645_/D sky130_fd_sc_hd__a2bb2o_4
X_19031_ _19029_/Y _19030_/X _18961_/X _19030_/X VGND VGND VPWR VPWR _23871_/D sky130_fd_sc_hd__a2bb2o_4
X_13455_ _13455_/A _19725_/A VGND VGND VPWR VPWR _13457_/B sky130_fd_sc_hd__or2_4
XFILLER_90_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19123__B1 _19056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12406_ _12406_/A VGND VGND VPWR VPWR _12407_/B sky130_fd_sc_hd__inv_2
XFILLER_16_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16174_ _14555_/B _16174_/B VGND VGND VPWR VPWR _16175_/D sky130_fd_sc_hd__and2_4
X_13386_ _13386_/A _13386_/B _13386_/C VGND VGND VPWR VPWR _13390_/B sky130_fd_sc_hd__and3_4
XFILLER_86_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15125_ _15125_/A VGND VGND VPWR VPWR _15125_/Y sky130_fd_sc_hd__inv_2
X_12337_ _24825_/Q VGND VGND VPWR VPWR _12337_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15056_ _14884_/Y _15190_/A _15022_/X _15055_/X VGND VGND VPWR VPWR _15057_/A sky130_fd_sc_hd__o22a_4
X_19933_ _19933_/A VGND VGND VPWR VPWR _22246_/B sky130_fd_sc_hd__inv_2
X_12268_ _25448_/Q _12255_/Y _12278_/C _24739_/Q VGND VGND VPWR VPWR _12271_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15160__B2 _24570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14007_ _14001_/A VGND VGND VPWR VPWR _14007_/X sky130_fd_sc_hd__buf_2
XANTENNA__17437__B1 _16720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22430__B1 _12318_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19864_ _19863_/Y _19859_/X _19841_/X _19859_/A VGND VGND VPWR VPWR _19864_/X sky130_fd_sc_hd__a2bb2o_4
X_12199_ _12199_/A VGND VGND VPWR VPWR _12199_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24965__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18815_ _18682_/A _18818_/B _18707_/X VGND VGND VPWR VPWR _18815_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__23246__A _23246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19795_ _19792_/Y _19793_/X _19794_/X _19793_/X VGND VGND VPWR VPWR _19795_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22150__A _15077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15074__A1_N _15073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18746_ _18656_/Y _18745_/X VGND VGND VPWR VPWR _18747_/A sky130_fd_sc_hd__or2_4
XFILLER_37_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15958_ _12257_/Y _15954_/X _15957_/X _15954_/X VGND VGND VPWR VPWR _24755_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14909_ _14908_/X _16855_/A _14908_/X _16855_/A VGND VGND VPWR VPWR _14909_/X sky130_fd_sc_hd__a2bb2o_4
X_18677_ _18677_/A VGND VGND VPWR VPWR _18680_/A sky130_fd_sc_hd__inv_2
X_15889_ _15886_/X _15887_/X _15739_/X _24788_/Q _15888_/X VGND VGND VPWR VPWR _15889_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12388__A _12179_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17628_ _17630_/B VGND VGND VPWR VPWR _17628_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23289__A2 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17559_ _17559_/A _17600_/C VGND VGND VPWR VPWR _17584_/C sky130_fd_sc_hd__or2_4
XANTENNA__19362__B1 _19294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20570_ _23939_/Q _18876_/X VGND VGND VPWR VPWR _20570_/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19229_ _13303_/B VGND VGND VPWR VPWR _19229_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22240_ _18291_/X _22236_/X _22239_/X VGND VGND VPWR VPWR _22240_/X sky130_fd_sc_hd__or3_4
XFILLER_69_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17125__C1 _17056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12201__A2 _22853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22325__A _17717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22171_ _22170_/X VGND VGND VPWR VPWR _22171_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21122_ _15662_/A _15662_/B _14406_/A _13813_/B VGND VGND VPWR VPWR _21335_/A sky130_fd_sc_hd__or4_4
XANTENNA__17428__B1 _16782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21053_ _21053_/A _15658_/A VGND VGND VPWR VPWR _21053_/X sky130_fd_sc_hd__and2_4
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20004_ _20004_/A VGND VGND VPWR VPWR _22243_/B sky130_fd_sc_hd__inv_2
XFILLER_101_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22060__A _22055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24635__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24812_ _24836_/CLK _24812_/D HRESETn VGND VGND VPWR VPWR _12345_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18928__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22724__A1 _24416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24743_ _25385_/CLK _24743_/D HRESETn VGND VGND VPWR VPWR _24743_/Q sky130_fd_sc_hd__dfrtp_4
X_21955_ _18261_/A _21953_/X _21954_/X _23336_/A _21636_/X VGND VGND VPWR VPWR _21955_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_28_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ _20905_/Y _20901_/Y VGND VGND VPWR VPWR _20906_/X sky130_fd_sc_hd__and2_4
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24674_ _24606_/CLK _16153_/X HRESETn VGND VGND VPWR VPWR _22183_/A sky130_fd_sc_hd__dfrtp_4
X_21886_ _21886_/A _21886_/B VGND VGND VPWR VPWR _21889_/B sky130_fd_sc_hd__or2_4
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21404__A _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23625_ _23598_/CLK _23625_/D VGND VGND VPWR VPWR _13325_/B sky130_fd_sc_hd__dfxtp_4
X_20837_ _24034_/Q VGND VGND VPWR VPWR _20837_/Y sky130_fd_sc_hd__inv_2
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14965__B2 _14900_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25494__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_246_0_HCLK clkbuf_8_247_0_HCLK/A VGND VGND VPWR VPWR _24427_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23556_ _23623_/CLK _23556_/D VGND VGND VPWR VPWR _19929_/A sky130_fd_sc_hd__dfxtp_4
X_20768_ _13120_/B _20761_/X _20767_/X VGND VGND VPWR VPWR _20768_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22507_ _22507_/A _22613_/B VGND VGND VPWR VPWR _22507_/Y sky130_fd_sc_hd__nor2_4
XFILLER_122_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25423__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12561__A2_N _12559_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23487_ _23453_/CLK _20119_/X VGND VGND VPWR VPWR _20117_/A sky130_fd_sc_hd__dfxtp_4
X_20699_ _20699_/A VGND VGND VPWR VPWR _20699_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18713__A _18705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ _13387_/A _13240_/B VGND VGND VPWR VPWR _13240_/X sky130_fd_sc_hd__or2_4
X_25226_ _23967_/CLK _25226_/D HRESETn VGND VGND VPWR VPWR _14001_/A sky130_fd_sc_hd__dfrtp_4
X_22438_ _17350_/B _22424_/A _12202_/A _22763_/A VGND VGND VPWR VPWR _22438_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13171_ _13190_/A _13171_/B VGND VGND VPWR VPWR _13171_/X sky130_fd_sc_hd__or2_4
X_25157_ _24102_/CLK _25157_/D HRESETn VGND VGND VPWR VPWR _23344_/B sky130_fd_sc_hd__dfrtp_4
X_22369_ _21624_/A _22367_/X _22368_/X VGND VGND VPWR VPWR _22369_/X sky130_fd_sc_hd__and3_4
XANTENNA__12761__A _25355_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12122_ _12166_/A _12119_/X _11862_/X _12119_/X VGND VGND VPWR VPWR _25457_/D sky130_fd_sc_hd__a2bb2o_4
X_24108_ _25205_/CLK _18890_/X HRESETn VGND VGND VPWR VPWR _24108_/Q sky130_fd_sc_hd__dfstp_4
X_25088_ _23978_/CLK _25088_/D HRESETn VGND VGND VPWR VPWR scl_oen_o_S4 sky130_fd_sc_hd__dfstp_4
XFILLER_85_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17419__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12053_ _12050_/X _15640_/B _15700_/C _13593_/D VGND VGND VPWR VPWR _12054_/A sky130_fd_sc_hd__or4_4
X_16930_ _16135_/Y _24257_/Q _16135_/Y _24257_/Q VGND VGND VPWR VPWR _16930_/X sky130_fd_sc_hd__a2bb2o_4
X_24039_ _24041_/CLK _24039_/D HRESETn VGND VGND VPWR VPWR _24039_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_5_9_0_HCLK_A clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16861_ _16861_/A VGND VGND VPWR VPWR _19780_/A sky130_fd_sc_hd__buf_2
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24376__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18600_ _16541_/Y _18599_/X _16541_/Y _24144_/Q VGND VGND VPWR VPWR _18600_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15812_ _15809_/A VGND VGND VPWR VPWR _15812_/X sky130_fd_sc_hd__buf_2
X_19580_ _22385_/A VGND VGND VPWR VPWR _19580_/Y sky130_fd_sc_hd__inv_2
X_16792_ _16792_/A VGND VGND VPWR VPWR _16792_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24305__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22715__A1 _24749_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22715__B2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18531_ _18464_/D _18523_/B VGND VGND VPWR VPWR _18532_/B sky130_fd_sc_hd__or2_4
X_12955_ _12955_/A _12955_/B VGND VGND VPWR VPWR _12956_/C sky130_fd_sc_hd__or2_4
X_15743_ HWDATA[15] VGND VGND VPWR VPWR _15743_/X sky130_fd_sc_hd__buf_2
X_11906_ _11872_/X _11905_/X _11896_/X _11904_/A VGND VGND VPWR VPWR _25503_/D sky130_fd_sc_hd__a22oi_4
X_18462_ _24160_/Q VGND VGND VPWR VPWR _18464_/C sky130_fd_sc_hd__inv_2
X_12886_ _12886_/A _12852_/X _12600_/X VGND VGND VPWR VPWR _12886_/X sky130_fd_sc_hd__or3_4
X_15674_ _16373_/A VGND VGND VPWR VPWR _15674_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_56_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15748__A3 _15747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17413_ _17413_/A VGND VGND VPWR VPWR _21355_/A sky130_fd_sc_hd__buf_2
XFILLER_61_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21314__A _21314_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11837_ HWDATA[6] VGND VGND VPWR VPWR _11838_/A sky130_fd_sc_hd__buf_2
X_14625_ _14624_/X VGND VGND VPWR VPWR _14625_/Y sky130_fd_sc_hd__inv_2
X_18393_ _18393_/A VGND VGND VPWR VPWR _18393_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12936__A _12936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19344__B1 _19232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16408__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11840__A _25512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14556_ _14555_/X VGND VGND VPWR VPWR _14586_/A sky130_fd_sc_hd__inv_2
X_17344_ _17344_/A VGND VGND VPWR VPWR _17370_/A sky130_fd_sc_hd__buf_2
XANTENNA__16158__B1 _15471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11768_ _11777_/A VGND VGND VPWR VPWR _11768_/X sky130_fd_sc_hd__buf_2
XANTENNA__21151__B1 _21314_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23940__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ _13497_/Y VGND VGND VPWR VPWR _13507_/X sky130_fd_sc_hd__buf_2
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14487_ _25103_/Q VGND VGND VPWR VPWR _14487_/Y sky130_fd_sc_hd__inv_2
X_17275_ _17277_/B VGND VGND VPWR VPWR _17276_/B sky130_fd_sc_hd__inv_2
XANTENNA__15905__B1 _15627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11699_ _11690_/X _11699_/B _11695_/X _11699_/D VGND VGND VPWR VPWR _11699_/X sky130_fd_sc_hd__or4_4
X_19014_ _19014_/A _19014_/B _19013_/X VGND VGND VPWR VPWR _19014_/X sky130_fd_sc_hd__or3_4
X_13438_ _13301_/X _13436_/X _13437_/X VGND VGND VPWR VPWR _13438_/X sky130_fd_sc_hd__and3_4
X_16226_ _16223_/Y _16225_/X _11796_/X _16225_/X VGND VGND VPWR VPWR _16226_/X sky130_fd_sc_hd__a2bb2o_4
X_16157_ _16087_/A VGND VGND VPWR VPWR _16157_/X sky130_fd_sc_hd__buf_2
X_13369_ _17452_/B _13369_/B VGND VGND VPWR VPWR _13369_/X sky130_fd_sc_hd__or2_4
XANTENNA__17239__A _17239_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16143__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15108_ _15322_/A VGND VGND VPWR VPWR _15309_/C sky130_fd_sc_hd__inv_2
X_16088_ _16088_/A VGND VGND VPWR VPWR _16088_/X sky130_fd_sc_hd__buf_2
XFILLER_88_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15039_ _15239_/A _24445_/Q _15239_/A _24445_/Q VGND VGND VPWR VPWR _15039_/X sky130_fd_sc_hd__a2bb2o_4
X_19916_ _19923_/A VGND VGND VPWR VPWR _19916_/X sky130_fd_sc_hd__buf_2
XFILLER_138_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22403__B1 _24710_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14892__B1 _15187_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19847_ _19859_/A VGND VGND VPWR VPWR _19847_/X sky130_fd_sc_hd__buf_2
XFILLER_64_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19778_ _19773_/Y _19776_/X _19777_/X _19776_/X VGND VGND VPWR VPWR _23612_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21208__B _21138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24046__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18729_ _18728_/X VGND VGND VPWR VPWR _18729_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16940__A1_N _16156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13007__A _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21740_ _21581_/X _21738_/X _21105_/A _21739_/X VGND VGND VPWR VPWR _21741_/B sky130_fd_sc_hd__o22a_4
XFILLER_92_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17702__A _17702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16397__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21671_ _21671_/A _21671_/B _21671_/C VGND VGND VPWR VPWR _21671_/X sky130_fd_sc_hd__and3_4
XFILLER_75_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19335__B1 _19313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23410_ _24209_/CLK _20323_/X VGND VGND VPWR VPWR _21978_/B sky130_fd_sc_hd__dfxtp_4
X_20622_ _15467_/Y _20605_/X _20619_/X _20621_/X VGND VGND VPWR VPWR _20623_/A sky130_fd_sc_hd__a211o_4
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24390_ _24356_/CLK _17058_/Y HRESETn VGND VGND VPWR VPWR _17022_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_127_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23341_ _24211_/Q _21979_/X _23339_/X _23340_/Y VGND VGND VPWR VPWR _23341_/X sky130_fd_sc_hd__a211o_4
X_20553_ _18874_/B _20552_/Y _20558_/C VGND VGND VPWR VPWR _20553_/X sky130_fd_sc_hd__and3_4
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_13_0_HCLK clkbuf_7_6_0_HCLK/X VGND VGND VPWR VPWR _23494_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_76_0_HCLK clkbuf_8_77_0_HCLK/A VGND VGND VPWR VPWR _24943_/CLK sky130_fd_sc_hd__clkbuf_1
X_23272_ _24802_/Q _23304_/B VGND VGND VPWR VPWR _23272_/X sky130_fd_sc_hd__or2_4
X_20484_ _20469_/A VGND VGND VPWR VPWR _20488_/B sky130_fd_sc_hd__buf_2
X_25011_ _25016_/CLK _15230_/Y HRESETn VGND VGND VPWR VPWR _25011_/Q sky130_fd_sc_hd__dfrtp_4
X_22223_ _13551_/Y _22727_/B _21162_/X VGND VGND VPWR VPWR _22223_/X sky130_fd_sc_hd__a21o_4
XFILLER_69_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18310__A1 _21658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24887__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22154_ _22154_/A _22298_/B VGND VGND VPWR VPWR _22154_/X sky130_fd_sc_hd__or2_4
XFILLER_69_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16321__B1 _15964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24816__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21105_ _21105_/A VGND VGND VPWR VPWR _22988_/A sky130_fd_sc_hd__buf_2
XANTENNA__23198__B2 _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19364__A _16781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22085_ _14991_/A _21073_/B _21326_/X VGND VGND VPWR VPWR _22085_/X sky130_fd_sc_hd__o21a_4
XFILLER_120_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22945__B2 _22280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21036_ _22835_/A VGND VGND VPWR VPWR _22664_/B sky130_fd_sc_hd__buf_2
XFILLER_134_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22987_ _23054_/A _22987_/B VGND VGND VPWR VPWR _22987_/Y sky130_fd_sc_hd__nor2_4
XFILLER_28_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15534__A1_N _15533_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22173__A2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12740_ _24767_/Q VGND VGND VPWR VPWR _12740_/Y sky130_fd_sc_hd__inv_2
X_21938_ _21458_/A _21938_/B VGND VGND VPWR VPWR _21938_/X sky130_fd_sc_hd__or2_4
XFILLER_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24726_ _24712_/CLK _16018_/X HRESETn VGND VGND VPWR VPWR _24726_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12671_ _12686_/A _12669_/X _12671_/C VGND VGND VPWR VPWR _25409_/D sky130_fd_sc_hd__and3_4
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24657_ _24517_/CLK _16208_/X HRESETn VGND VGND VPWR VPWR _16207_/A sky130_fd_sc_hd__dfrtp_4
X_21869_ _24739_/Q _21025_/A _15854_/X _24811_/Q _15544_/X VGND VGND VPWR VPWR _21869_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_70_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16228__A _11800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19326__B1 _19212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12756__A _25381_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ HWDATA[7] VGND VGND VPWR VPWR _16057_/A sky130_fd_sc_hd__buf_2
XFILLER_42_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23608_ _23453_/CLK _19791_/X VGND VGND VPWR VPWR _19789_/A sky130_fd_sc_hd__dfxtp_4
X_15390_ _15390_/A _15409_/A VGND VGND VPWR VPWR _15390_/X sky130_fd_sc_hd__or2_4
XFILLER_70_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21133__B1 _13467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24588_ _24984_/CLK _24588_/D HRESETn VGND VGND VPWR VPWR _15089_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _14340_/X VGND VGND VPWR VPWR _14341_/Y sky130_fd_sc_hd__inv_2
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21684__A1 _13795_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23539_ _23394_/CLK _23539_/D VGND VGND VPWR VPWR _19977_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22881__B1 _22797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21684__B2 _18261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17060_ _17060_/A _17060_/B VGND VGND VPWR VPWR _17061_/A sky130_fd_sc_hd__or2_4
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14272_ _21548_/A _14271_/X _13803_/X _14271_/X VGND VGND VPWR VPWR _14272_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16011_ _16009_/Y _16010_/X _11761_/X _16010_/X VGND VGND VPWR VPWR _24729_/D sky130_fd_sc_hd__a2bb2o_4
X_13223_ _13309_/A _13223_/B _13222_/X VGND VGND VPWR VPWR _13223_/X sky130_fd_sc_hd__and3_4
XANTENNA__21436__A1 _23314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25209_ _25093_/CLK _14138_/X HRESETn VGND VGND VPWR VPWR _14117_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__11801__A1_N _11798_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13154_ _13168_/A _13154_/B _13153_/X VGND VGND VPWR VPWR _13154_/X sky130_fd_sc_hd__and3_4
XFILLER_88_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16312__B1 _15955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24557__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12105_ _12104_/Y _12102_/X _11829_/X _12102_/X VGND VGND VPWR VPWR _12105_/X sky130_fd_sc_hd__a2bb2o_4
X_13085_ _12991_/B _13097_/B VGND VGND VPWR VPWR _13092_/B sky130_fd_sc_hd__or2_4
X_17962_ _17944_/X _17959_/X _18021_/A _24236_/Q _17960_/X VGND VGND VPWR VPWR _24236_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19701_ _19699_/Y _19697_/X _19700_/X _19697_/X VGND VGND VPWR VPWR _23638_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22412__B _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12036_ _12036_/A VGND VGND VPWR VPWR _12036_/Y sky130_fd_sc_hd__inv_2
X_16913_ _16906_/X _16908_/X _16913_/C _16913_/D VGND VGND VPWR VPWR _16913_/X sky130_fd_sc_hd__or4_4
XANTENNA__21309__A _16723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17893_ _17893_/A VGND VGND VPWR VPWR _17893_/Y sky130_fd_sc_hd__inv_2
X_19632_ _19632_/A VGND VGND VPWR VPWR _19632_/X sky130_fd_sc_hd__buf_2
XANTENNA__11835__A _25513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16844_ _16840_/A VGND VGND VPWR VPWR _16844_/X sky130_fd_sc_hd__buf_2
XFILLER_120_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19563_ _22342_/B _19562_/X _11930_/X _19562_/X VGND VGND VPWR VPWR _19563_/X sky130_fd_sc_hd__a2bb2o_4
X_16775_ _15008_/Y _16773_/X _16604_/X _16773_/X VGND VGND VPWR VPWR _16775_/X sky130_fd_sc_hd__a2bb2o_4
X_13987_ _14042_/A VGND VGND VPWR VPWR _14012_/A sky130_fd_sc_hd__buf_2
XFILLER_111_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18514_ _18517_/A _18514_/B _18514_/C VGND VGND VPWR VPWR _24169_/D sky130_fd_sc_hd__and3_4
XFILLER_0_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15726_ _15548_/X _15713_/X _15725_/X _24867_/Q _15711_/X VGND VGND VPWR VPWR _15726_/X
+ sky130_fd_sc_hd__a32o_4
X_12938_ _12937_/X VGND VGND VPWR VPWR _12938_/Y sky130_fd_sc_hd__inv_2
X_19494_ _19494_/A VGND VGND VPWR VPWR _19494_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16379__B1 _16285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23243__B _23069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21911__A2 _21910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18429__A1_N _16237_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18445_ _16261_/Y _24148_/Q _21322_/A _18475_/C VGND VGND VPWR VPWR _18445_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15657_ _21074_/B VGND VGND VPWR VPWR _15658_/A sky130_fd_sc_hd__buf_2
XANTENNA__25345__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12869_ _12840_/Y _12856_/X VGND VGND VPWR VPWR _12869_/X sky130_fd_sc_hd__or2_4
XANTENNA__25181__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14608_ _14561_/A _14560_/X VGND VGND VPWR VPWR _14608_/Y sky130_fd_sc_hd__nand2_4
X_18376_ _24183_/Q VGND VGND VPWR VPWR _18376_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21124__B1 _14182_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15588_ _15588_/A VGND VGND VPWR VPWR _15588_/X sky130_fd_sc_hd__buf_2
XANTENNA__20883__A _20900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12385__B _12385_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17327_ _17253_/Y _17320_/B _17279_/X _17324_/Y VGND VGND VPWR VPWR _17327_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17879__B1 _16955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14539_ _14539_/A VGND VGND VPWR VPWR _14539_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17258_ _17236_/Y _17258_/B VGND VGND VPWR VPWR _17282_/B sky130_fd_sc_hd__or2_4
XFILLER_128_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16209_ _23004_/A VGND VGND VPWR VPWR _16209_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22624__B1 _24854_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17189_ _17188_/Y VGND VGND VPWR VPWR _17349_/A sky130_fd_sc_hd__buf_2
XFILLER_115_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24980__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24298__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24227__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17416__B _14223_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23137__C _23136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22910_ _17254_/C _22908_/X _12778_/A _22909_/X VGND VGND VPWR VPWR _22910_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23890_ _25488_/CLK _23890_/D VGND VGND VPWR VPWR _23890_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16082__A2 _15668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22841_ _12228_/Y _22268_/X _16728_/A _12341_/Y _22840_/X VGND VGND VPWR VPWR _22842_/B
+ sky130_fd_sc_hd__o32a_4
XANTENNA__22155__A2 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19556__B1 _19462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22772_ _22770_/X _22771_/X _22479_/X _16033_/A _22480_/X VGND VGND VPWR VPWR _22772_/X
+ sky130_fd_sc_hd__a32o_4
X_24511_ _24541_/CLK _24511_/D HRESETn VGND VGND VPWR VPWR _24511_/Q sky130_fd_sc_hd__dfrtp_4
X_21723_ _21556_/X _21723_/B VGND VGND VPWR VPWR _21723_/X sky130_fd_sc_hd__and2_4
XANTENNA__25086__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25491_ _23711_/CLK _25491_/D HRESETn VGND VGND VPWR VPWR _19995_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19308__B1 _19307_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24442_ _25002_/CLK _16774_/X HRESETn VGND VGND VPWR VPWR _15013_/A sky130_fd_sc_hd__dfrtp_4
X_21654_ _21456_/A _21654_/B VGND VGND VPWR VPWR _21654_/X sky130_fd_sc_hd__or2_4
XANTENNA__25015__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21115__B1 _21106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20605_ _20604_/Y VGND VGND VPWR VPWR _20605_/X sky130_fd_sc_hd__buf_2
X_24373_ _24373_/CLK _24373_/D HRESETn VGND VGND VPWR VPWR _17036_/A sky130_fd_sc_hd__dfrtp_4
X_21585_ _21581_/X _21582_/X _22280_/A _21584_/X VGND VGND VPWR VPWR _21586_/B sky130_fd_sc_hd__o22a_4
XFILLER_138_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23324_ _24565_/Q _23166_/X _21326_/X VGND VGND VPWR VPWR _23324_/X sky130_fd_sc_hd__o21a_4
X_20536_ _20536_/A VGND VGND VPWR VPWR _23931_/D sky130_fd_sc_hd__inv_2
XFILLER_138_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23255_ _23255_/A VGND VGND VPWR VPWR _23255_/Y sky130_fd_sc_hd__inv_2
X_20467_ _20467_/A _20474_/B _20481_/C VGND VGND VPWR VPWR _20468_/A sky130_fd_sc_hd__or3_4
X_22206_ _22193_/X _19088_/Y VGND VGND VPWR VPWR _22206_/X sky130_fd_sc_hd__or2_4
XANTENNA__22091__A1 _24539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23186_ _23185_/X VGND VGND VPWR VPWR _23186_/Y sky130_fd_sc_hd__inv_2
X_20398_ _20231_/C _17462_/Y _19219_/X VGND VGND VPWR VPWR _20399_/A sky130_fd_sc_hd__or3_4
XANTENNA__24650__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22137_ _16352_/A _22654_/A VGND VGND VPWR VPWR _22137_/X sky130_fd_sc_hd__or2_4
XFILLER_133_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22068_ _22068_/A _22068_/B VGND VGND VPWR VPWR _22069_/C sky130_fd_sc_hd__or2_4
XFILLER_59_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12867__C1 _12866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19795__B1 _19794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18598__B2 _18789_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13910_ _13909_/X VGND VGND VPWR VPWR _13918_/C sky130_fd_sc_hd__inv_2
X_21019_ _21019_/A VGND VGND VPWR VPWR _22929_/A sky130_fd_sc_hd__buf_2
X_14890_ _14890_/A VGND VGND VPWR VPWR _14890_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13841_ _13543_/Y _13839_/X _13840_/X _13839_/X VGND VGND VPWR VPWR _25247_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_121_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_243_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13772_ _13771_/X VGND VGND VPWR VPWR _16725_/A sky130_fd_sc_hd__buf_2
X_16560_ _16560_/A VGND VGND VPWR VPWR _16560_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15511_ _15490_/X VGND VGND VPWR VPWR _15511_/X sky130_fd_sc_hd__buf_2
X_12723_ _12704_/B VGND VGND VPWR VPWR _12724_/B sky130_fd_sc_hd__inv_2
XFILLER_91_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24709_ _24356_/CLK _16062_/X HRESETn VGND VGND VPWR VPWR _24709_/Q sky130_fd_sc_hd__dfrtp_4
X_16491_ _16474_/A VGND VGND VPWR VPWR _16491_/X sky130_fd_sc_hd__buf_2
XFILLER_71_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18230_ _18230_/A _18230_/B VGND VGND VPWR VPWR _18231_/A sky130_fd_sc_hd__or2_4
X_12654_ _12517_/Y _12652_/X _12653_/X VGND VGND VPWR VPWR _12654_/Y sky130_fd_sc_hd__a21oi_4
X_15442_ _14280_/X _20525_/A _15441_/Y _13957_/B _15438_/X VGND VGND VPWR VPWR _24959_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21799__A _21469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18161_ _18097_/A _18161_/B _18160_/X VGND VGND VPWR VPWR _18161_/X sky130_fd_sc_hd__and3_4
XANTENNA__15797__A _15817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _12524_/Y _24868_/Q _25408_/Q _12584_/Y VGND VGND VPWR VPWR _12589_/C sky130_fd_sc_hd__a2bb2o_4
X_15373_ _15373_/A VGND VGND VPWR VPWR _15373_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15012__D _15012_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17112_ _17108_/A _17105_/X _17112_/C VGND VGND VPWR VPWR _17112_/X sky130_fd_sc_hd__and3_4
XANTENNA__22407__B _22407_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14324_ _14329_/A _23344_/B _25156_/Q VGND VGND VPWR VPWR _25157_/D sky130_fd_sc_hd__a21o_4
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18092_ _17995_/A VGND VGND VPWR VPWR _18191_/A sky130_fd_sc_hd__buf_2
XANTENNA__21311__B _22927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24738__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14255_ _14255_/A VGND VGND VPWR VPWR _21139_/B sky130_fd_sc_hd__buf_2
X_17043_ _17043_/A VGND VGND VPWR VPWR _17043_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18901__A _18900_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13206_ _13345_/A _13206_/B VGND VGND VPWR VPWR _13206_/X sky130_fd_sc_hd__or2_4
X_14186_ _14185_/Y VGND VGND VPWR VPWR _20479_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24391__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13137_ _20804_/A _20799_/A _13137_/C _13136_/X VGND VGND VPWR VPWR _13137_/X sky130_fd_sc_hd__or4_4
XFILLER_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18994_ _18991_/Y _18989_/X _18993_/X _18989_/X VGND VGND VPWR VPWR _18994_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24320__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13068_ _12349_/Y _13052_/B _13010_/A _13065_/Y VGND VGND VPWR VPWR _13068_/X sky130_fd_sc_hd__a211o_4
X_17945_ _17929_/A _17945_/B VGND VGND VPWR VPWR _17945_/X sky130_fd_sc_hd__or2_4
X_12019_ _12019_/A _12019_/B VGND VGND VPWR VPWR _12021_/A sky130_fd_sc_hd__and2_4
XANTENNA__12322__B2 _12321_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17876_ _17876_/A VGND VGND VPWR VPWR _17876_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19615_ _19615_/A VGND VGND VPWR VPWR _19615_/X sky130_fd_sc_hd__buf_2
X_16827_ _24416_/Q VGND VGND VPWR VPWR _16827_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25526__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17252__A _17252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23334__B2 _13598_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19546_ _23689_/Q VGND VGND VPWR VPWR _19546_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16758_ _16733_/A VGND VGND VPWR VPWR _16773_/A sky130_fd_sc_hd__buf_2
XFILLER_0_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15709_ _15709_/A _15703_/A VGND VGND VPWR VPWR _15740_/A sky130_fd_sc_hd__or2_4
X_19477_ _22020_/B _19471_/X _11939_/X _19476_/X VGND VGND VPWR VPWR _23714_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16689_ _16687_/Y _16683_/X _15747_/X _16688_/X VGND VGND VPWR VPWR _24479_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15024__B1 _25005_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_26_0_HCLK clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18428_ _21322_/A _18475_/C _22089_/A _18427_/Y VGND VGND VPWR VPWR _18428_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16772__B1 _11821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18359_ _18359_/A VGND VGND VPWR VPWR _18359_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22845__B1 _12559_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18083__A _18221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21370_ _14620_/D _18270_/X _17700_/C VGND VGND VPWR VPWR _21370_/X sky130_fd_sc_hd__o21a_4
XANTENNA__20118__A _20105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24479__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20321_ _20320_/X VGND VGND VPWR VPWR _20326_/A sky130_fd_sc_hd__buf_2
XFILLER_134_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24408__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23040_ _21295_/X VGND VGND VPWR VPWR _23040_/X sky130_fd_sc_hd__buf_2
X_20252_ _19844_/X _19084_/D _19845_/C VGND VGND VPWR VPWR _20252_/X sky130_fd_sc_hd__or3_4
XFILLER_115_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23270__B1 _24837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22333__A _21942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12561__B2 _24847_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20183_ _20181_/Y _20182_/X _20096_/X _20182_/X VGND VGND VPWR VPWR _20183_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24061__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24991_ _24984_/CLK _24991_/D HRESETn VGND VGND VPWR VPWR _24991_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13510__B1 _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19642__A _19642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23942_ _25122_/CLK _23942_/D HRESETn VGND VGND VPWR VPWR _23942_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25267__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23873_ _23689_/CLK _19026_/X VGND VGND VPWR VPWR _23873_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22824_ _22824_/A VGND VGND VPWR VPWR _22824_/X sky130_fd_sc_hd__buf_2
XANTENNA__12077__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17500__A1_N _25517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22755_ _12927_/A _22753_/X _22754_/X VGND VGND VPWR VPWR _22755_/X sky130_fd_sc_hd__o21a_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21706_ _21704_/X _21706_/B _21048_/B VGND VGND VPWR VPWR _21706_/X sky130_fd_sc_hd__or3_4
XANTENNA__23089__B1 _12539_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25474_ _24376_/CLK _12062_/X HRESETn VGND VGND VPWR VPWR _23344_/A sky130_fd_sc_hd__dfrtp_4
X_22686_ _22786_/A _22682_/X _23056_/A _22685_/X VGND VGND VPWR VPWR _22687_/A sky130_fd_sc_hd__o22a_4
XANTENNA__13577__B1 _13575_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21412__A _21069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24425_ _24457_/CLK _24425_/D HRESETn VGND VGND VPWR VPWR _14919_/A sky130_fd_sc_hd__dfrtp_4
X_21637_ _21200_/B VGND VGND VPWR VPWR _21995_/A sky130_fd_sc_hd__buf_2
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21639__B2 _22390_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22300__A2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12370_ _25344_/Q _12368_/Y _12990_/B _24827_/Q VGND VGND VPWR VPWR _12371_/D sky130_fd_sc_hd__a2bb2o_4
X_24356_ _24356_/CLK _24356_/D HRESETn VGND VGND VPWR VPWR _24356_/Q sky130_fd_sc_hd__dfrtp_4
X_21568_ _21567_/X VGND VGND VPWR VPWR _21568_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24831__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23307_ _24630_/Q _21519_/B VGND VGND VPWR VPWR _23307_/X sky130_fd_sc_hd__or2_4
X_20519_ _20519_/A _20519_/B VGND VGND VPWR VPWR _20519_/X sky130_fd_sc_hd__or2_4
XFILLER_125_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24287_ _24285_/CLK _17675_/X HRESETn VGND VGND VPWR VPWR _17517_/A sky130_fd_sc_hd__dfrtp_4
X_21499_ _21496_/X _21499_/B _21498_/X VGND VGND VPWR VPWR _21499_/X sky130_fd_sc_hd__and3_4
XFILLER_5_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24149__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_46_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_93_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_14040_ _13989_/X _14039_/Y _14040_/C _14040_/D VGND VGND VPWR VPWR _14041_/A sky130_fd_sc_hd__or4_4
XFILLER_88_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12472__C _12282_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23238_ _24429_/Q _22135_/X _22797_/X _23237_/X VGND VGND VPWR VPWR _23239_/C sky130_fd_sc_hd__a211o_4
XANTENNA__23261__B1 _12328_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17337__A _17249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23169_ _23133_/A _23169_/B _23169_/C VGND VGND VPWR VPWR _23169_/X sky130_fd_sc_hd__and3_4
XFILLER_121_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14829__B1 _14226_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15991_ _15991_/A _15991_/B _15991_/C _15991_/D VGND VGND VPWR VPWR _15992_/B sky130_fd_sc_hd__or4_4
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12304__B2 _24823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17730_ _17729_/Y VGND VGND VPWR VPWR _17730_/X sky130_fd_sc_hd__buf_2
X_14942_ _25000_/Q VGND VGND VPWR VPWR _14942_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20698__A _20676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17661_ _17557_/Y _17577_/Y VGND VGND VPWR VPWR _17695_/A sky130_fd_sc_hd__or2_4
XFILLER_75_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14873_ _14869_/Y _14872_/Y _14864_/X VGND VGND VPWR VPWR _14873_/X sky130_fd_sc_hd__o21a_4
XFILLER_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19400_ _19400_/A VGND VGND VPWR VPWR _19401_/A sky130_fd_sc_hd__inv_2
XFILLER_21_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22119__A2 _22083_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23316__A1 _25451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16612_ _16611_/Y _16609_/X _16528_/X _16609_/X VGND VGND VPWR VPWR _24507_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13824_ _13562_/Y _13822_/X _11804_/X _13822_/X VGND VGND VPWR VPWR _25256_/D sky130_fd_sc_hd__a2bb2o_4
X_17592_ _17591_/X VGND VGND VPWR VPWR _24308_/D sky130_fd_sc_hd__inv_2
XFILLER_47_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21327__B1 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19331_ _17933_/B VGND VGND VPWR VPWR _19331_/Y sky130_fd_sc_hd__inv_2
X_16543_ _16795_/A _16459_/B VGND VGND VPWR VPWR _16550_/A sky130_fd_sc_hd__nor2_4
X_13755_ _13755_/A _13752_/X _20043_/A _14697_/A VGND VGND VPWR VPWR _20077_/A sky130_fd_sc_hd__or4_4
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12706_ _12706_/A _12706_/B VGND VGND VPWR VPWR _12707_/B sky130_fd_sc_hd__or2_4
X_19262_ _23788_/Q VGND VGND VPWR VPWR _19262_/Y sky130_fd_sc_hd__inv_2
X_16474_ _16474_/A VGND VGND VPWR VPWR _16474_/X sky130_fd_sc_hd__buf_2
X_13686_ _11663_/Y _13685_/X VGND VGND VPWR VPWR _13686_/X sky130_fd_sc_hd__or2_4
XANTENNA__16754__B1 _16405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24919__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18213_ _18181_/A _18213_/B _18213_/C VGND VGND VPWR VPWR _18217_/B sky130_fd_sc_hd__and3_4
X_15425_ _15425_/A VGND VGND VPWR VPWR _15425_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21322__A _21322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12637_ _12657_/A _12635_/X _12637_/C VGND VGND VPWR VPWR _25417_/D sky130_fd_sc_hd__and3_4
X_19193_ _19193_/A VGND VGND VPWR VPWR _19193_/Y sky130_fd_sc_hd__inv_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23240__C _23235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22137__B _22654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18144_ _18176_/A _18144_/B _18144_/C VGND VGND VPWR VPWR _18145_/C sky130_fd_sc_hd__and3_4
X_12568_ _12567_/Y _24856_/Q _12567_/Y _24856_/Q VGND VGND VPWR VPWR _12568_/X sky130_fd_sc_hd__a2bb2o_4
X_15356_ _15356_/A _15354_/A VGND VGND VPWR VPWR _15357_/C sky130_fd_sc_hd__or2_4
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24572__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14307_ _14296_/B VGND VGND VPWR VPWR _14307_/X sky130_fd_sc_hd__buf_2
XFILLER_7_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18075_ _18175_/A _23889_/Q VGND VGND VPWR VPWR _18076_/C sky130_fd_sc_hd__or2_4
X_12499_ _12499_/A _12499_/B VGND VGND VPWR VPWR _12499_/X sky130_fd_sc_hd__or2_4
X_15287_ _24995_/Q _15315_/A VGND VGND VPWR VPWR _15287_/X sky130_fd_sc_hd__or2_4
XFILLER_32_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24501__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17026_ _17026_/A VGND VGND VPWR VPWR _17026_/Y sky130_fd_sc_hd__inv_2
X_14238_ _14238_/A VGND VGND VPWR VPWR _14238_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22153__A _23170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14169_ _25119_/Q VGND VGND VPWR VPWR _14169_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16151__A _22183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_3_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_113_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18977_ _16786_/X VGND VGND VPWR VPWR _18977_/X sky130_fd_sc_hd__buf_2
XFILLER_100_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15493__B1 HADDR[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15990__A _24734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17928_ _17928_/A VGND VGND VPWR VPWR _17928_/X sky130_fd_sc_hd__buf_2
XANTENNA__19462__A _19055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17859_ _17846_/X _17850_/X VGND VGND VPWR VPWR _17862_/B sky130_fd_sc_hd__or2_4
XFILLER_27_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25360__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20870_ _13663_/B VGND VGND VPWR VPWR _20870_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21318__B1 _22885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19529_ _19527_/Y _19528_/X _11952_/X _19528_/X VGND VGND VPWR VPWR _19529_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21869__A1 _24739_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11806__B1 _11804_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18734__A1 _18675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22540_ _22540_/A VGND VGND VPWR VPWR _23226_/B sky130_fd_sc_hd__buf_2
XFILLER_34_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22328__A _21944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22471_ _23035_/A VGND VGND VPWR VPWR _22472_/B sky130_fd_sc_hd__buf_2
XFILLER_37_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24210_ _25508_/CLK _18266_/X HRESETn VGND VGND VPWR VPWR _18265_/A sky130_fd_sc_hd__dfrtp_4
X_21422_ _21043_/Y VGND VGND VPWR VPWR _21422_/X sky130_fd_sc_hd__buf_2
X_25190_ _25172_/CLK _14215_/X HRESETn VGND VGND VPWR VPWR _14214_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_135_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24141_ _24133_/CLK _18716_/Y HRESETn VGND VGND VPWR VPWR _24141_/Q sky130_fd_sc_hd__dfrtp_4
X_21353_ _14876_/Y _21352_/X _14238_/Y _14221_/A VGND VGND VPWR VPWR _21359_/B sky130_fd_sc_hd__o22a_4
XANTENNA__24242__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20304_ _20298_/Y VGND VGND VPWR VPWR _20304_/X sky130_fd_sc_hd__buf_2
X_24072_ _24069_/CLK _24072_/D HRESETn VGND VGND VPWR VPWR _20515_/B sky130_fd_sc_hd__dfrtp_4
X_21284_ _21284_/A VGND VGND VPWR VPWR _21285_/A sky130_fd_sc_hd__buf_2
XFILLER_89_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23023_ _12259_/Y _22268_/X _22712_/X _12368_/Y _22840_/X VGND VGND VPWR VPWR _23024_/B
+ sky130_fd_sc_hd__o32a_4
X_20235_ _13214_/B VGND VGND VPWR VPWR _20235_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16061__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22998__A _22998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20166_ _20165_/Y _20161_/X _20123_/X _20161_/A VGND VGND VPWR VPWR _23469_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25448__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17307__D _17247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20097_ _20094_/Y _20095_/X _20096_/X _20095_/X VGND VGND VPWR VPWR _20097_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24974_ _24977_/CLK _15397_/X HRESETn VGND VGND VPWR VPWR _24974_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21407__A _21320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23925_ _24077_/CLK _20977_/X HRESETn VGND VGND VPWR VPWR _23925_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20311__A _20298_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15236__B1 _15199_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11870_ _11870_/A VGND VGND VPWR VPWR _11900_/A sky130_fd_sc_hd__inv_2
XFILLER_79_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25030__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23856_ _23854_/CLK _19074_/X VGND VGND VPWR VPWR _13337_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13798__B1 _13797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11652__B _11970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22807_ _22778_/X _22781_/X _22789_/Y _22806_/X VGND VGND VPWR VPWR HRDATA[16] sky130_fd_sc_hd__a211o_4
X_20999_ _23962_/Q _23963_/Q _21000_/B VGND VGND VPWR VPWR _20999_/X sky130_fd_sc_hd__o21a_4
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23787_ _24398_/CLK _19269_/X VGND VGND VPWR VPWR _19268_/A sky130_fd_sc_hd__dfxtp_4
X_13540_ _15677_/A _13540_/B VGND VGND VPWR VPWR _14619_/A sky130_fd_sc_hd__or2_4
XFILLER_129_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25526_ _25526_/CLK _11786_/X HRESETn VGND VGND VPWR VPWR _25526_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15539__B2 _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22738_ _21040_/A _22737_/X _22396_/C _24857_/Q _22547_/X VGND VGND VPWR VPWR _22738_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_40_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16538__A2_N _16461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13471_ _13471_/A VGND VGND VPWR VPWR _13471_/Y sky130_fd_sc_hd__inv_2
X_25457_ _24097_/CLK _25457_/D HRESETn VGND VGND VPWR VPWR _12121_/A sky130_fd_sc_hd__dfrtp_4
X_22669_ _22669_/A VGND VGND VPWR VPWR _22669_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12764__A _25373_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12422_ _12422_/A VGND VGND VPWR VPWR _12422_/Y sky130_fd_sc_hd__inv_2
X_15210_ _14961_/X _15210_/B _15210_/C VGND VGND VPWR VPWR _15211_/B sky130_fd_sc_hd__or3_4
XFILLER_40_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12222__B1 _12220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24408_ _24998_/CLK _24408_/D HRESETn VGND VGND VPWR VPWR _14922_/A sky130_fd_sc_hd__dfrtp_4
X_16190_ _16189_/Y _16187_/X _11746_/X _16187_/X VGND VGND VPWR VPWR _16190_/X sky130_fd_sc_hd__a2bb2o_4
X_25388_ _25400_/CLK _12739_/Y HRESETn VGND VGND VPWR VPWR _25388_/Q sky130_fd_sc_hd__dfrtp_4
X_12353_ _12352_/Y _24820_/Q _12352_/Y _24820_/Q VGND VGND VPWR VPWR _12353_/X sky130_fd_sc_hd__a2bb2o_4
X_15141_ _15134_/X _15141_/B _15138_/X _15140_/X VGND VGND VPWR VPWR _15162_/B sky130_fd_sc_hd__or4_4
XANTENNA__19547__A _15766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24339_ _24334_/CLK _24339_/D HRESETn VGND VGND VPWR VPWR _17240_/A sky130_fd_sc_hd__dfrtp_4
X_15072_ _15187_/A _15072_/B VGND VGND VPWR VPWR _15165_/A sky130_fd_sc_hd__or2_4
XANTENNA__13798__A1_N _23336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12284_ _12284_/A VGND VGND VPWR VPWR _12285_/C sky130_fd_sc_hd__inv_2
XFILLER_114_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23234__B1 _22834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23069__A _24558_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14023_ _14023_/A _14003_/B VGND VGND VPWR VPWR _14025_/C sky130_fd_sc_hd__or2_4
X_18900_ _13736_/X _19084_/D _19822_/C VGND VGND VPWR VPWR _18900_/X sky130_fd_sc_hd__or3_4
XANTENNA__17067__A _17384_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13722__B1 _13714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13595__A _13595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12525__B2 _24868_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19880_ _19880_/A VGND VGND VPWR VPWR _19880_/X sky130_fd_sc_hd__buf_2
X_18831_ _16533_/Y _18681_/A _16533_/Y _18681_/A VGND VGND VPWR VPWR _18831_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_133_0_HCLK clkbuf_7_66_0_HCLK/X VGND VGND VPWR VPWR _23905_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18661__B1 _16620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15475__B1 _15474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_196_0_HCLK clkbuf_7_98_0_HCLK/X VGND VGND VPWR VPWR _24893_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18762_ _18759_/A _18758_/B _18761_/X VGND VGND VPWR VPWR _18762_/X sky130_fd_sc_hd__and3_4
X_15974_ _15788_/X _15969_/X _11818_/A _24746_/Q _15933_/A VGND VGND VPWR VPWR _15974_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_27_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17713_ _17713_/A VGND VGND VPWR VPWR _17713_/X sky130_fd_sc_hd__buf_2
X_14925_ _25014_/Q VGND VGND VPWR VPWR _15067_/C sky130_fd_sc_hd__inv_2
X_18693_ _18693_/A _18693_/B VGND VGND VPWR VPWR _18693_/X sky130_fd_sc_hd__or2_4
XFILLER_29_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20220__B1 _19715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17644_ _17642_/A _17641_/B _17643_/Y VGND VGND VPWR VPWR _17644_/X sky130_fd_sc_hd__and3_4
X_14856_ _14828_/X _14855_/X _24944_/Q _14835_/X VGND VGND VPWR VPWR _14856_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__16975__B1 _16054_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13807_ _21366_/A _13804_/X _13515_/X _13804_/X VGND VGND VPWR VPWR _25259_/D sky130_fd_sc_hd__a2bb2o_4
X_17575_ _17662_/A _17662_/B _17574_/Y _17499_/Y VGND VGND VPWR VPWR _17575_/X sky130_fd_sc_hd__or4_4
X_14787_ _18177_/A VGND VGND VPWR VPWR _18017_/A sky130_fd_sc_hd__buf_2
X_11999_ _11991_/A _11991_/B _11998_/Y VGND VGND VPWR VPWR _12001_/A sky130_fd_sc_hd__o21a_4
XFILLER_44_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19314_ _19309_/Y _19312_/X _19313_/X _19312_/X VGND VGND VPWR VPWR _19314_/X sky130_fd_sc_hd__a2bb2o_4
X_16526_ _16523_/Y _16524_/X _16525_/X _16524_/X VGND VGND VPWR VPWR _16526_/X sky130_fd_sc_hd__a2bb2o_4
X_13738_ _13738_/A VGND VGND VPWR VPWR _13739_/B sky130_fd_sc_hd__inv_2
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24753__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19245_ _22354_/B _19244_/X _16863_/X _19244_/X VGND VGND VPWR VPWR _23796_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16457_ _24565_/Q VGND VGND VPWR VPWR _16457_/Y sky130_fd_sc_hd__inv_2
X_13669_ _13668_/X VGND VGND VPWR VPWR _13669_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12674__A _12567_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15408_ _15408_/A _15406_/Y _15407_/X VGND VGND VPWR VPWR _15408_/X sky130_fd_sc_hd__and3_4
XFILLER_34_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19176_ _19175_/Y VGND VGND VPWR VPWR _19176_/X sky130_fd_sc_hd__buf_2
X_16388_ _24593_/Q VGND VGND VPWR VPWR _16388_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18127_ _18191_/A _18127_/B _18126_/X VGND VGND VPWR VPWR _18127_/X sky130_fd_sc_hd__and3_4
X_15339_ _15315_/A VGND VGND VPWR VPWR _15339_/X sky130_fd_sc_hd__buf_2
X_18058_ _18058_/A _18058_/B _18057_/X VGND VGND VPWR VPWR _18058_/X sky130_fd_sc_hd__or3_4
XANTENNA__12300__A1_N _12299_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20039__B1 _19995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17009_ _24382_/Q VGND VGND VPWR VPWR _17048_/B sky130_fd_sc_hd__inv_2
XFILLER_132_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22579__A2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12516__B2 _12527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_92_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_92_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20020_ _20018_/Y _20014_/X _20019_/X _20014_/A VGND VGND VPWR VPWR _20020_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22611__A _22574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15466__B1 _14414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21971_ _18230_/A _21970_/X VGND VGND VPWR VPWR _21971_/Y sky130_fd_sc_hd__nand2_4
XFILLER_73_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11753__A _11753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20922_ _24053_/Q _20922_/B VGND VGND VPWR VPWR _20922_/Y sky130_fd_sc_hd__nor2_4
XFILLER_66_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23710_ _23398_/CLK _23710_/D VGND VGND VPWR VPWR _23710_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15769__A1 _15749_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24690_ _24692_/CLK _16111_/X HRESETn VGND VGND VPWR VPWR _24690_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20853_ _20851_/A _20847_/X _20852_/X VGND VGND VPWR VPWR _20853_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_54_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23641_ _23649_/CLK _19693_/X VGND VGND VPWR VPWR _13317_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22503__A2 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23572_ _23623_/CLK _23572_/D VGND VGND VPWR VPWR _19887_/A sky130_fd_sc_hd__dfxtp_4
X_20784_ _24021_/Q _20783_/B _20783_/Y VGND VGND VPWR VPWR _20784_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16718__B1 _16717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24494__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22523_ _22523_/A VGND VGND VPWR VPWR _22523_/X sky130_fd_sc_hd__buf_2
XANTENNA__19380__B2 _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25311_ _25309_/CLK _25311_/D HRESETn VGND VGND VPWR VPWR _25311_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16056__A _24710_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24423__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22454_ _22453_/X VGND VGND VPWR VPWR _22462_/B sky130_fd_sc_hd__inv_2
X_25242_ _25263_/CLK _25242_/D HRESETn VGND VGND VPWR VPWR _25242_/Q sky130_fd_sc_hd__dfrtp_4
X_21405_ _21369_/X _21370_/X _22505_/A _21404_/X VGND VGND VPWR VPWR _21405_/X sky130_fd_sc_hd__a211o_4
X_25173_ _24151_/CLK _14274_/X HRESETn VGND VGND VPWR VPWR _14273_/A sky130_fd_sc_hd__dfrtp_4
X_22385_ _22385_/A _22389_/B VGND VGND VPWR VPWR _22385_/X sky130_fd_sc_hd__or2_4
XFILLER_135_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24124_ _24117_/CLK _24124_/D HRESETn VGND VGND VPWR VPWR _18677_/A sky130_fd_sc_hd__dfrtp_4
X_21336_ _21336_/A VGND VGND VPWR VPWR _21351_/B sky130_fd_sc_hd__inv_2
XFILLER_68_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24055_ _24055_/CLK _24055_/D HRESETn VGND VGND VPWR VPWR _20931_/A sky130_fd_sc_hd__dfrtp_4
X_21267_ _13598_/C _18270_/X VGND VGND VPWR VPWR _21267_/Y sky130_fd_sc_hd__nor2_4
XFILLER_137_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23006_ _24524_/Q _22393_/X _15668_/A _23005_/X VGND VGND VPWR VPWR _23007_/C sky130_fd_sc_hd__a211o_4
X_20218_ _20216_/Y _20212_/X _19758_/X _20217_/X VGND VGND VPWR VPWR _20218_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18643__B1 _16592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25282__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21198_ _20335_/A _19582_/X VGND VGND VPWR VPWR _21198_/X sky130_fd_sc_hd__or2_4
XFILLER_132_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_206_0_HCLK clkbuf_8_207_0_HCLK/A VGND VGND VPWR VPWR _24811_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__14451__A1_N _14182_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20149_ _20161_/A VGND VGND VPWR VPWR _20149_/X sky130_fd_sc_hd__buf_2
XFILLER_106_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25211__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12971_ _12845_/B _12970_/X VGND VGND VPWR VPWR _12975_/B sky130_fd_sc_hd__or2_4
X_24957_ _24957_/CLK _15445_/X HRESETn VGND VGND VPWR VPWR _24957_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14710_ _14676_/A VGND VGND VPWR VPWR _14710_/Y sky130_fd_sc_hd__inv_2
X_11922_ _11922_/A VGND VGND VPWR VPWR _19612_/A sky130_fd_sc_hd__buf_2
XFILLER_131_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23908_ _23905_/CLK _23908_/D VGND VGND VPWR VPWR _23908_/Q sky130_fd_sc_hd__dfxtp_4
X_15690_ _15687_/B _15687_/C VGND VGND VPWR VPWR _15690_/X sky130_fd_sc_hd__or2_4
XFILLER_73_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24888_ _24889_/CLK _24888_/D HRESETn VGND VGND VPWR VPWR _24888_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14641_ _17957_/A _14641_/B _14638_/X _18006_/A VGND VGND VPWR VPWR _14641_/X sky130_fd_sc_hd__and4_4
X_11853_ _16359_/A VGND VGND VPWR VPWR _11853_/X sky130_fd_sc_hd__buf_2
X_23839_ _25488_/CLK _23839_/D VGND VGND VPWR VPWR _19119_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_82_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17350__A _17350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17360_ _17196_/A _17359_/Y VGND VGND VPWR VPWR _17360_/X sky130_fd_sc_hd__or2_4
X_11784_ HWDATA[19] VGND VGND VPWR VPWR _11784_/X sky130_fd_sc_hd__buf_2
X_14572_ _14572_/A _14571_/Y VGND VGND VPWR VPWR _14573_/A sky130_fd_sc_hd__or2_4
XFILLER_92_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21702__B1 _24706_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16311_ _16288_/X VGND VGND VPWR VPWR _16311_/X sky130_fd_sc_hd__buf_2
X_13523_ _25170_/Q _13522_/X VGND VGND VPWR VPWR _13524_/B sky130_fd_sc_hd__or2_4
X_25509_ _25508_/CLK _11859_/X HRESETn VGND VGND VPWR VPWR _25509_/Q sky130_fd_sc_hd__dfrtp_4
X_17291_ _17222_/Y _17256_/X _17346_/B VGND VGND VPWR VPWR _17291_/X sky130_fd_sc_hd__or3_4
XANTENNA__24164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19030_ _19030_/A VGND VGND VPWR VPWR _19030_/X sky130_fd_sc_hd__buf_2
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16242_ _11818_/A VGND VGND VPWR VPWR _16242_/X sky130_fd_sc_hd__buf_2
XFILLER_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13454_ _13454_/A _13454_/B _13453_/X VGND VGND VPWR VPWR _13454_/X sky130_fd_sc_hd__or3_4
XFILLER_51_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15301__C _15073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12405_ _12290_/X _13008_/B VGND VGND VPWR VPWR _12406_/A sky130_fd_sc_hd__or2_4
X_13385_ _13417_/A _19696_/A VGND VGND VPWR VPWR _13386_/C sky130_fd_sc_hd__or2_4
X_16173_ _16173_/A _16173_/B VGND VGND VPWR VPWR _16174_/B sky130_fd_sc_hd__and2_4
XFILLER_126_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15124_ _24980_/Q _15122_/Y _15390_/A _15126_/A VGND VGND VPWR VPWR _15124_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12336_ _25340_/Q VGND VGND VPWR VPWR _13054_/A sky130_fd_sc_hd__inv_2
XFILLER_31_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11838__A _11838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_16_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_12267_ _12266_/Y _24765_/Q _12266_/Y _24765_/Q VGND VGND VPWR VPWR _12271_/B sky130_fd_sc_hd__a2bb2o_4
X_15055_ _15055_/A _15055_/B _15055_/C _15054_/X VGND VGND VPWR VPWR _15055_/X sky130_fd_sc_hd__or4_4
X_19932_ _19929_/Y _19931_/X _19612_/X _19931_/X VGND VGND VPWR VPWR _23556_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14006_ _14006_/A _14006_/B _25221_/Q _14005_/Y VGND VGND VPWR VPWR _14006_/X sky130_fd_sc_hd__and4_4
X_19863_ _23581_/Q VGND VGND VPWR VPWR _19863_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18634__B1 _16618_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22430__A1 _12204_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12198_ _12198_/A _12198_/B _12195_/X _12198_/D VGND VGND VPWR VPWR _12198_/X sky130_fd_sc_hd__or4_4
XANTENNA__22430__B2 _21529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18814_ _18682_/B _18820_/B VGND VGND VPWR VPWR _18818_/B sky130_fd_sc_hd__or2_4
XANTENNA__17525__A _24295_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19794_ _16879_/A VGND VGND VPWR VPWR _19794_/X sky130_fd_sc_hd__buf_2
XANTENNA__23246__B _21017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22150__B _22927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18745_ _18691_/X _18756_/B VGND VGND VPWR VPWR _18745_/X sky130_fd_sc_hd__or2_4
XFILLER_114_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21047__A _21306_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15957_ HWDATA[20] VGND VGND VPWR VPWR _15957_/X sky130_fd_sc_hd__buf_2
XFILLER_62_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14908_ _15061_/D VGND VGND VPWR VPWR _14908_/X sky130_fd_sc_hd__buf_2
XANTENNA__19740__A _18254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18676_ _18674_/Y _18675_/X VGND VGND VPWR VPWR _18676_/X sky130_fd_sc_hd__or2_4
X_15888_ _15863_/A VGND VGND VPWR VPWR _15888_/X sky130_fd_sc_hd__buf_2
XANTENNA__24934__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17627_ _17541_/Y _17626_/X VGND VGND VPWR VPWR _17630_/B sky130_fd_sc_hd__or2_4
X_14839_ _14838_/X VGND VGND VPWR VPWR _14839_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14884__A pwm_S6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17260__A _17260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17558_ _17557_/Y VGND VGND VPWR VPWR _17611_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_5_26_0_HCLK_A clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16509_ _16508_/Y _16504_/X _16238_/X _16504_/X VGND VGND VPWR VPWR _16509_/X sky130_fd_sc_hd__a2bb2o_4
X_17489_ _17489_/A _17489_/B _17485_/X _17488_/X VGND VGND VPWR VPWR _17489_/X sky130_fd_sc_hd__or4_4
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19228_ _19226_/Y _19222_/X _19136_/X _19227_/X VGND VGND VPWR VPWR _23802_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19159_ _19159_/A VGND VGND VPWR VPWR _19159_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20802__A1_N _20680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16604__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16540__A1_N _16539_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22170_ _21560_/X _22168_/X _21566_/X _22169_/X VGND VGND VPWR VPWR _22170_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12851__B _12799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21121_ _23921_/Q VGND VGND VPWR VPWR _21121_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21052_ _15665_/A VGND VGND VPWR VPWR _21729_/A sky130_fd_sc_hd__buf_2
XANTENNA__15639__A2_N _15563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20003_ _22333_/B _20002_/X _19975_/X _20002_/X VGND VGND VPWR VPWR _20003_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24811_ _24811_/CLK _15837_/X HRESETn VGND VGND VPWR VPWR _24811_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22185__B1 _21103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_36_0_HCLK clkbuf_8_37_0_HCLK/A VGND VGND VPWR VPWR _25264_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__19050__B1 _18977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24742_ _25385_/CLK _15980_/X HRESETn VGND VGND VPWR VPWR _22400_/A sky130_fd_sc_hd__dfrtp_4
X_21954_ _19546_/Y _21995_/A VGND VGND VPWR VPWR _21954_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_99_0_HCLK clkbuf_8_99_0_HCLK/A VGND VGND VPWR VPWR _24318_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21932__B1 _18298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24675__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23172__A _22798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20905_ _24049_/Q VGND VGND VPWR VPWR _20905_/Y sky130_fd_sc_hd__inv_2
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ _21398_/A VGND VGND VPWR VPWR _21885_/X sky130_fd_sc_hd__buf_2
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24673_ _24673_/CLK _16155_/X HRESETn VGND VGND VPWR VPWR _22144_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_43_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24604__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _20814_/X VGND VGND VPWR VPWR _20836_/X sky130_fd_sc_hd__buf_2
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23624_ _23598_/CLK _19741_/X VGND VGND VPWR VPWR _13360_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20767_ _20767_/A _20767_/B VGND VGND VPWR VPWR _20767_/X sky130_fd_sc_hd__and2_4
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23555_ _23623_/CLK _19934_/X VGND VGND VPWR VPWR _19933_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22506_ _13831_/Y _22506_/B VGND VGND VPWR VPWR _22506_/X sky130_fd_sc_hd__and2_4
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23486_ _23478_/CLK _20121_/X VGND VGND VPWR VPWR _23486_/Q sky130_fd_sc_hd__dfxtp_4
X_20698_ _20676_/X VGND VGND VPWR VPWR _20698_/X sky130_fd_sc_hd__buf_2
XFILLER_109_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22437_ _22963_/A VGND VGND VPWR VPWR _22763_/A sky130_fd_sc_hd__buf_2
X_25225_ _23967_/CLK _25225_/D HRESETn VGND VGND VPWR VPWR _13989_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13170_ _18344_/A _13170_/B VGND VGND VPWR VPWR _13172_/B sky130_fd_sc_hd__or2_4
X_22368_ _21618_/A _22368_/B VGND VGND VPWR VPWR _22368_/X sky130_fd_sc_hd__or2_4
X_25156_ _25205_/CLK _14328_/X HRESETn VGND VGND VPWR VPWR _25156_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20036__A _20036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25463__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12121_ _12121_/A VGND VGND VPWR VPWR _12166_/A sky130_fd_sc_hd__inv_2
X_21319_ _14944_/A _21312_/X _22997_/A _21318_/X VGND VGND VPWR VPWR _21320_/C sky130_fd_sc_hd__a211o_4
X_24107_ _25205_/CLK _18891_/X HRESETn VGND VGND VPWR VPWR _24107_/Q sky130_fd_sc_hd__dfstp_4
X_25087_ _24322_/CLK _25087_/D HRESETn VGND VGND VPWR VPWR sda_oen_o_S4 sky130_fd_sc_hd__dfstp_4
X_22299_ _24440_/Q _21293_/X _22885_/A VGND VGND VPWR VPWR _22299_/X sky130_fd_sc_hd__o21a_4
X_12052_ _12052_/A _12052_/B VGND VGND VPWR VPWR _13593_/D sky130_fd_sc_hd__or2_4
X_24038_ _24581_/CLK _20859_/Y HRESETn VGND VGND VPWR VPWR _24038_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22889__C _22889_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16860_ _16858_/Y _16859_/X RsRx_S0 _16859_/X VGND VGND VPWR VPWR _16860_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15811_ _12366_/Y _15809_/X _11781_/X _15809_/X VGND VGND VPWR VPWR _15811_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16791_ _16790_/Y _16730_/A _16717_/X _16730_/A VGND VGND VPWR VPWR _24434_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18530_ _18530_/A VGND VGND VPWR VPWR _18530_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22715__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15742_ _15742_/A VGND VGND VPWR VPWR _15742_/X sky130_fd_sc_hd__buf_2
XANTENNA__19041__B1 _19018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12954_ _12954_/A _12953_/Y VGND VGND VPWR VPWR _12956_/B sky130_fd_sc_hd__or2_4
XFILLER_133_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11905_ _11896_/X _11899_/Y _11904_/Y VGND VGND VPWR VPWR _11905_/X sky130_fd_sc_hd__o21a_4
X_18461_ _18461_/A VGND VGND VPWR VPWR _18461_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15673_ _22884_/B VGND VGND VPWR VPWR _16373_/A sky130_fd_sc_hd__buf_2
X_12885_ _12884_/X VGND VGND VPWR VPWR _25381_/D sky130_fd_sc_hd__inv_2
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24345__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_7_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17412_ _14807_/A VGND VGND VPWR VPWR _20662_/A sky130_fd_sc_hd__buf_2
X_14624_ _14613_/A _13637_/A _14623_/X VGND VGND VPWR VPWR _14624_/X sky130_fd_sc_hd__a21o_4
X_11836_ _11794_/X VGND VGND VPWR VPWR _11836_/X sky130_fd_sc_hd__buf_2
X_18392_ _16179_/Y _24176_/Q _16179_/Y _24176_/Q VGND VGND VPWR VPWR _18392_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21314__B _21314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17343_ _17342_/X VGND VGND VPWR VPWR _17343_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14555_ _13769_/Y _14555_/B VGND VGND VPWR VPWR _14555_/X sky130_fd_sc_hd__or2_4
X_11767_ HWDATA[24] VGND VGND VPWR VPWR _11767_/X sky130_fd_sc_hd__buf_2
XANTENNA__21151__A1 _16539_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _13505_/Y _13501_/X _11842_/X _13501_/X VGND VGND VPWR VPWR _25299_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17274_ _17261_/B _17260_/X VGND VGND VPWR VPWR _17277_/B sky130_fd_sc_hd__or2_4
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14486_ _21708_/A _14481_/X _14403_/X _14481_/X VGND VGND VPWR VPWR _14486_/X sky130_fd_sc_hd__a2bb2o_4
X_11698_ _13693_/C _24226_/Q _13702_/A _11697_/Y VGND VGND VPWR VPWR _11699_/D sky130_fd_sc_hd__o22a_4
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22426__A _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19013_ _13617_/Y _13613_/X _14659_/A VGND VGND VPWR VPWR _19013_/X sky130_fd_sc_hd__or3_4
X_16225_ _16225_/A VGND VGND VPWR VPWR _16225_/X sky130_fd_sc_hd__buf_2
XANTENNA__21330__A _14377_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13437_ _13270_/A _23437_/Q VGND VGND VPWR VPWR _13437_/X sky130_fd_sc_hd__or2_4
XFILLER_31_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18644__A1_N _16587_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23980__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16156_ _24672_/Q VGND VGND VPWR VPWR _16156_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13368_ _13198_/X _13367_/X _25316_/Q _13258_/X VGND VGND VPWR VPWR _25316_/D sky130_fd_sc_hd__o22a_4
X_15107_ _15097_/X _15100_/X _15107_/C _15106_/X VGND VGND VPWR VPWR _15121_/C sky130_fd_sc_hd__or4_4
X_12319_ _25330_/Q _24815_/Q _12991_/B _12318_/Y VGND VGND VPWR VPWR _12319_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19735__A _19729_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16087_ _16087_/A VGND VGND VPWR VPWR _16088_/A sky130_fd_sc_hd__buf_2
XANTENNA__25133__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13299_ _13402_/A _23841_/Q VGND VGND VPWR VPWR _13299_/X sky130_fd_sc_hd__or2_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15038_ _14947_/Y VGND VGND VPWR VPWR _15239_/A sky130_fd_sc_hd__buf_2
X_19915_ _19915_/A VGND VGND VPWR VPWR _22076_/B sky130_fd_sc_hd__inv_2
XANTENNA__22403__A1 _22271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18659__A1_N _24524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22403__B2 _21067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17255__A _22659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19846_ _19846_/A VGND VGND VPWR VPWR _19859_/A sky130_fd_sc_hd__inv_2
XFILLER_122_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16999__A2_N _17036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16989_ _16989_/A _16989_/B _16989_/C _16988_/X VGND VGND VPWR VPWR _16990_/D sky130_fd_sc_hd__or4_4
X_19777_ _19777_/A VGND VGND VPWR VPWR _19777_/X sky130_fd_sc_hd__buf_2
XFILLER_3_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12399__A _12399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_252_0_HCLK clkbuf_7_126_0_HCLK/X VGND VGND VPWR VPWR _24457_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15841__B1 _15840_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18728_ _18675_/X _18728_/B VGND VGND VPWR VPWR _18728_/X sky130_fd_sc_hd__or2_4
XFILLER_64_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18659_ _24524_/Q _18658_/Y _16572_/Y _24133_/Q VGND VGND VPWR VPWR _18660_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24086__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21670_ _21670_/A _19990_/Y VGND VGND VPWR VPWR _21671_/C sky130_fd_sc_hd__or2_4
XANTENNA__24015__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20621_ _20621_/A _20621_/B _20611_/C VGND VGND VPWR VPWR _20621_/X sky130_fd_sc_hd__and3_4
XFILLER_51_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18814__A _18682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23340_ _18259_/Y _23340_/B VGND VGND VPWR VPWR _23340_/Y sky130_fd_sc_hd__nor2_4
X_20552_ _18873_/A _18873_/B VGND VGND VPWR VPWR _20552_/Y sky130_fd_sc_hd__nand2_4
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23271_ _23271_/A _23271_/B VGND VGND VPWR VPWR _23281_/B sky130_fd_sc_hd__and2_4
X_20483_ _20519_/A _20483_/B VGND VGND VPWR VPWR _24073_/D sky130_fd_sc_hd__or2_4
XFILLER_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12862__A _12600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22222_ _22222_/A VGND VGND VPWR VPWR _22222_/Y sky130_fd_sc_hd__inv_2
X_25010_ _25010_/CLK _25010_/D HRESETn VGND VGND VPWR VPWR _15233_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18846__B1 _16485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22153_ _23170_/A _22153_/B _22153_/C VGND VGND VPWR VPWR _22153_/X sky130_fd_sc_hd__and3_4
XANTENNA__20756__A1_N _20743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19645__A _18996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21104_ _15551_/B VGND VGND VPWR VPWR _21105_/A sky130_fd_sc_hd__buf_2
XFILLER_82_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23198__A2 _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22084_ _15126_/A _23082_/B VGND VGND VPWR VPWR _22087_/B sky130_fd_sc_hd__or2_4
XFILLER_47_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_62_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21035_ _21030_/X _21034_/Y _12980_/A _21030_/X VGND VGND VPWR VPWR _21035_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22945__A2 _22824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24856__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14939__D _14938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15832__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12102__A _12119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22986_ _22783_/X _22984_/X _22786_/X _22985_/X VGND VGND VPWR VPWR _22987_/B sky130_fd_sc_hd__o22a_4
XFILLER_76_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24725_ _24712_/CLK _16020_/X HRESETn VGND VGND VPWR VPWR _24725_/Q sky130_fd_sc_hd__dfrtp_4
X_21937_ _17717_/A _21937_/B VGND VGND VPWR VPWR _21937_/X sky130_fd_sc_hd__or2_4
XFILLER_83_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12670_ _12670_/A _12670_/B VGND VGND VPWR VPWR _12671_/C sky130_fd_sc_hd__or2_4
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24656_ _24654_/CLK _16210_/X HRESETn VGND VGND VPWR VPWR _23004_/A sky130_fd_sc_hd__dfrtp_4
X_21868_ _16156_/Y _21418_/X _22644_/B _11844_/Y _21570_/X VGND VGND VPWR VPWR _21868_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_54_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ _23478_/CLK _19795_/X VGND VGND VPWR VPWR _19792_/A sky130_fd_sc_hd__dfxtp_4
X_20819_ _16719_/Y _20815_/X _21209_/A _20818_/X VGND VGND VPWR VPWR _20819_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21133__A1 _13517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21799_ _21469_/A _21799_/B _21799_/C VGND VGND VPWR VPWR _21799_/X sky130_fd_sc_hd__or3_4
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24587_ _24984_/CLK _24587_/D HRESETn VGND VGND VPWR VPWR _15147_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ _14337_/Y _14338_/Y _14339_/Y _14336_/C VGND VGND VPWR VPWR _14340_/X sky130_fd_sc_hd__or4_4
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22881__A1 _24520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23538_ _23682_/CLK _19983_/X VGND VGND VPWR VPWR _23538_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21150__A _16448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15899__B1 _15756_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14271_ _14271_/A VGND VGND VPWR VPWR _14271_/X sky130_fd_sc_hd__buf_2
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23469_ _23581_/CLK _23469_/D VGND VGND VPWR VPWR _20165_/A sky130_fd_sc_hd__dfxtp_4
X_16010_ _16002_/X VGND VGND VPWR VPWR _16010_/X sky130_fd_sc_hd__buf_2
X_13222_ _13270_/A _13222_/B VGND VGND VPWR VPWR _13222_/X sky130_fd_sc_hd__or2_4
XFILLER_104_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25208_ _25122_/CLK _25208_/D HRESETn VGND VGND VPWR VPWR _14117_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18837__B1 _16535_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13153_ _13180_/A _23644_/Q VGND VGND VPWR VPWR _13153_/X sky130_fd_sc_hd__or2_4
X_25139_ _24945_/CLK _25139_/D HRESETn VGND VGND VPWR VPWR _14386_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_124_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12104_ _25464_/Q VGND VGND VPWR VPWR _12104_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13084_ _13096_/A _13084_/B VGND VGND VPWR VPWR _13097_/B sky130_fd_sc_hd__or2_4
X_17961_ _17960_/X VGND VGND VPWR VPWR _18021_/A sky130_fd_sc_hd__inv_2
XANTENNA__15088__A1_N _24973_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14874__A1 _14868_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22397__B1 _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12035_ _12033_/Y _12029_/X _12036_/A _12034_/X VGND VGND VPWR VPWR _12035_/X sky130_fd_sc_hd__a2bb2o_4
X_16912_ _22395_/A _24252_/Q _16149_/Y _16911_/Y VGND VGND VPWR VPWR _16913_/D sky130_fd_sc_hd__o22a_4
X_19700_ _19055_/X VGND VGND VPWR VPWR _19700_/X sky130_fd_sc_hd__buf_2
XANTENNA__17075__A _17384_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17892_ _17900_/A _17889_/X _24243_/Q _17891_/Y VGND VGND VPWR VPWR _17904_/A sky130_fd_sc_hd__o22a_4
XFILLER_120_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16076__B1 _15480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24597__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16843_ _14922_/Y _16840_/X _16521_/X _16840_/X VGND VGND VPWR VPWR _24408_/D sky130_fd_sc_hd__a2bb2o_4
X_19631_ _19631_/A VGND VGND VPWR VPWR _19631_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15823__B1 _24819_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24526__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19562_ _19574_/A VGND VGND VPWR VPWR _19562_/X sky130_fd_sc_hd__buf_2
XFILLER_24_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16774_ _15013_/Y _16770_/X _16600_/X _16773_/X VGND VGND VPWR VPWR _16774_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13986_ _14003_/B VGND VGND VPWR VPWR _13995_/A sky130_fd_sc_hd__inv_2
XFILLER_59_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18513_ _18460_/B _18517_/B VGND VGND VPWR VPWR _18514_/C sky130_fd_sc_hd__nand2_4
X_15725_ HWDATA[25] VGND VGND VPWR VPWR _15725_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19565__B2 _19562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12937_ _12799_/X _12931_/X _12884_/A _12933_/Y VGND VGND VPWR VPWR _12937_/X sky130_fd_sc_hd__a211o_4
X_19493_ _20338_/A _18278_/D _19492_/X VGND VGND VPWR VPWR _19494_/A sky130_fd_sc_hd__or3_4
XANTENNA__23243__C _23005_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12947__A _12842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_82_0_HCLK clkbuf_8_83_0_HCLK/A VGND VGND VPWR VPWR _25043_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__11851__A HWDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18444_ _18444_/A _18439_/X _18444_/C _18444_/D VGND VGND VPWR VPWR _18444_/X sky130_fd_sc_hd__or4_4
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15656_ _15653_/A VGND VGND VPWR VPWR _21074_/B sky130_fd_sc_hd__buf_2
X_12868_ _12868_/A VGND VGND VPWR VPWR _25385_/D sky130_fd_sc_hd__inv_2
XFILLER_18_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14607_ _14563_/B _14606_/Y _14599_/X _14602_/X _13573_/A VGND VGND VPWR VPWR _25073_/D
+ sky130_fd_sc_hd__a32o_4
X_11819_ _11815_/Y _11816_/X _11818_/X _11816_/X VGND VGND VPWR VPWR _25518_/D sky130_fd_sc_hd__a2bb2o_4
X_18375_ _18374_/Y _18372_/X _24183_/Q _18372_/X VGND VGND VPWR VPWR _18375_/X sky130_fd_sc_hd__a2bb2o_4
X_15587_ _15587_/A VGND VGND VPWR VPWR _15587_/Y sky130_fd_sc_hd__inv_2
X_12799_ _12799_/A VGND VGND VPWR VPWR _12799_/X sky130_fd_sc_hd__buf_2
XFILLER_14_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21124__B2 _21352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12385__C _12266_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17326_ _17306_/X _17321_/X _17325_/X VGND VGND VPWR VPWR _24345_/D sky130_fd_sc_hd__and3_4
XFILLER_18_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14538_ _14041_/Y _14043_/Y _14538_/C _14538_/D VGND VGND VPWR VPWR _14539_/A sky130_fd_sc_hd__or4_4
XANTENNA__25385__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_2_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__16000__B1 _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17257_ _17257_/A _17222_/Y _17239_/X _17256_/X VGND VGND VPWR VPWR _17258_/B sky130_fd_sc_hd__or4_4
XANTENNA__13778__A _11733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14469_ HWDATA[1] VGND VGND VPWR VPWR _14470_/A sky130_fd_sc_hd__buf_2
XANTENNA__25314__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16208_ _16207_/Y _16205_/X _11771_/X _16205_/X VGND VGND VPWR VPWR _16208_/X sky130_fd_sc_hd__a2bb2o_4
X_17188_ _24335_/Q VGND VGND VPWR VPWR _17188_/Y sky130_fd_sc_hd__inv_2
X_16139_ _16137_/Y _16138_/X _11818_/X _16138_/X VGND VGND VPWR VPWR _16139_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18598__A1_N _16594_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21060__B1 _21050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19829_ _19836_/A VGND VGND VPWR VPWR _19829_/X sky130_fd_sc_hd__buf_2
XFILLER_69_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24267__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15814__B1 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16082__A3 _15927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22840_ _21863_/X VGND VGND VPWR VPWR _22840_/X sky130_fd_sc_hd__buf_2
X_22771_ _24615_/Q _22626_/B VGND VGND VPWR VPWR _22771_/X sky130_fd_sc_hd__or2_4
XANTENNA__12857__A _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11761__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24510_ _24553_/CLK _24510_/D HRESETn VGND VGND VPWR VPWR _16603_/A sky130_fd_sc_hd__dfrtp_4
X_21722_ _16261_/Y _16449_/A _24570_/Q _16723_/A VGND VGND VPWR VPWR _21723_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25490_ _23388_/CLK _11956_/X HRESETn VGND VGND VPWR VPWR _19885_/A sky130_fd_sc_hd__dfrtp_4
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21653_ _21649_/X _21652_/X _17722_/X VGND VGND VPWR VPWR _21661_/B sky130_fd_sc_hd__o21a_4
XFILLER_80_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24441_ _24998_/CLK _16775_/X HRESETn VGND VGND VPWR VPWR _24441_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20604_ _17403_/A VGND VGND VPWR VPWR _20604_/Y sky130_fd_sc_hd__inv_2
X_21584_ _21584_/A _21019_/A VGND VGND VPWR VPWR _21584_/X sky130_fd_sc_hd__and2_4
XANTENNA__12800__B1 _12799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24372_ _24364_/CLK _24372_/D HRESETn VGND VGND VPWR VPWR _24372_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20535_ _14169_/Y _20533_/X _14452_/X _20534_/X VGND VGND VPWR VPWR _20536_/A sky130_fd_sc_hd__a211o_4
XFILLER_138_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23323_ _23323_/A _22832_/B VGND VGND VPWR VPWR _23323_/X sky130_fd_sc_hd__or2_4
XANTENNA__25055__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16064__A _16528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20466_ _13851_/A _20466_/B _13853_/A VGND VGND VPWR VPWR _20481_/C sky130_fd_sc_hd__or3_4
X_23254_ _21409_/A _23252_/X _22826_/X _23253_/X VGND VGND VPWR VPWR _23255_/A sky130_fd_sc_hd__o22a_4
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22205_ _22200_/A _22205_/B VGND VGND VPWR VPWR _22207_/B sky130_fd_sc_hd__or2_4
XANTENNA__22091__A2 _21026_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23185_ _23106_/X _23184_/X _23040_/X _24730_/Q _22972_/X VGND VGND VPWR VPWR _23185_/X
+ sky130_fd_sc_hd__a32o_4
X_20397_ _23378_/Q VGND VGND VPWR VPWR _20397_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22513__B _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12513__A2_N _24873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22136_ _21525_/A VGND VGND VPWR VPWR _22654_/A sky130_fd_sc_hd__buf_2
XFILLER_47_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22067_ _14682_/B _20258_/Y VGND VGND VPWR VPWR _22067_/X sky130_fd_sc_hd__or2_4
XFILLER_59_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16058__B1 _16057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24690__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21018_ _21018_/A VGND VGND VPWR VPWR _21019_/A sky130_fd_sc_hd__buf_2
XANTENNA__20968__B _14380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13840_ _11842_/A VGND VGND VPWR VPWR _13840_/X sky130_fd_sc_hd__buf_2
XANTENNA__23344__B _23344_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13771_ _24936_/Q VGND VGND VPWR VPWR _13771_/X sky130_fd_sc_hd__buf_2
XANTENNA__15820__A3 _11800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12767__A _25363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22969_ _22470_/X _22967_/X _22968_/X _12526_/A _22766_/X VGND VGND VPWR VPWR _22970_/B
+ sky130_fd_sc_hd__a32o_4
X_15510_ _11729_/D VGND VGND VPWR VPWR _15510_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_69_0_HCLK clkbuf_7_69_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_69_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12722_ _12706_/B _12720_/Y _12721_/X VGND VGND VPWR VPWR _25394_/D sky130_fd_sc_hd__and3_4
XFILLER_15_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24708_ _24356_/CLK _16065_/X HRESETn VGND VGND VPWR VPWR _24708_/Q sky130_fd_sc_hd__dfrtp_4
X_16490_ _16490_/A VGND VGND VPWR VPWR _16490_/Y sky130_fd_sc_hd__inv_2
X_15441_ _15441_/A _15434_/X VGND VGND VPWR VPWR _15441_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__23360__A _21003_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23919__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12653_ _12631_/B VGND VGND VPWR VPWR _12653_/X sky130_fd_sc_hd__buf_2
XFILLER_54_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24639_ _24162_/CLK _24639_/D HRESETn VGND VGND VPWR VPWR _22089_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18160_ _18058_/A _18160_/B _18159_/X VGND VGND VPWR VPWR _18160_/X sky130_fd_sc_hd__or3_4
XFILLER_19_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ _15372_/A _15369_/B _15371_/Y VGND VGND VPWR VPWR _24979_/D sky130_fd_sc_hd__and3_4
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _24862_/Q VGND VGND VPWR VPWR _12584_/Y sky130_fd_sc_hd__inv_2
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17111_ _17105_/A _17105_/B VGND VGND VPWR VPWR _17112_/C sky130_fd_sc_hd__nand2_4
XFILLER_129_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ _25158_/Q _13644_/X _14307_/X _25304_/Q _14305_/Y VGND VGND VPWR VPWR _25158_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13598__A _11710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18091_ _18220_/A _18089_/X _18090_/X VGND VGND VPWR VPWR _18096_/B sky130_fd_sc_hd__and3_4
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17042_ _24364_/Q VGND VGND VPWR VPWR _17044_/B sky130_fd_sc_hd__inv_2
X_14254_ _14254_/A VGND VGND VPWR VPWR _14254_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13205_ _13212_/A VGND VGND VPWR VPWR _13345_/A sky130_fd_sc_hd__buf_2
XFILLER_109_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14185_ _20493_/A VGND VGND VPWR VPWR _14185_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24778__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13136_ _13136_/A _24021_/Q _13118_/X _20783_/B VGND VGND VPWR VPWR _13136_/X sky130_fd_sc_hd__or4_4
XFILLER_97_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18993_ _19642_/A VGND VGND VPWR VPWR _18993_/X sky130_fd_sc_hd__buf_2
XANTENNA__24707__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15318__A _15318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11846__A _15766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13067_ _13049_/A _13067_/B _13066_/X VGND VGND VPWR VPWR _13067_/X sky130_fd_sc_hd__and3_4
X_17944_ _17928_/X _17944_/B _17943_/X VGND VGND VPWR VPWR _17944_/X sky130_fd_sc_hd__or3_4
XFILLER_61_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14222__A _14195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12018_ _12014_/Y _12017_/X _12014_/Y _12017_/X VGND VGND VPWR VPWR _12018_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17875_ _17747_/C _17848_/X _17790_/A _17872_/Y VGND VGND VPWR VPWR _17876_/A sky130_fd_sc_hd__a211o_4
XFILLER_61_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24360__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19614_ _23667_/Q VGND VGND VPWR VPWR _19614_/Y sky130_fd_sc_hd__inv_2
X_16826_ _16823_/Y _16825_/X _15739_/X _16825_/X VGND VGND VPWR VPWR _16826_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16757_ _15030_/Y _16753_/X _16410_/X _16753_/X VGND VGND VPWR VPWR _24450_/D sky130_fd_sc_hd__a2bb2o_4
X_19545_ _19543_/Y _19539_/X _19407_/X _19544_/X VGND VGND VPWR VPWR _19545_/X sky130_fd_sc_hd__a2bb2o_4
X_13969_ _13969_/A _13905_/X VGND VGND VPWR VPWR _13970_/C sky130_fd_sc_hd__and2_4
XANTENNA__17549__B1 _11850_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16969__A1_N _24724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21345__B2 _16453_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15708_ _15708_/A VGND VGND VPWR VPWR _15709_/A sky130_fd_sc_hd__buf_2
XFILLER_111_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16688_ _16664_/A VGND VGND VPWR VPWR _16688_/X sky130_fd_sc_hd__buf_2
X_19476_ _19470_/Y VGND VGND VPWR VPWR _19476_/X sky130_fd_sc_hd__buf_2
XFILLER_62_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15639_ _15638_/Y _15563_/A _15480_/X _15563_/A VGND VGND VPWR VPWR _24880_/D sky130_fd_sc_hd__a2bb2o_4
X_18427_ _18581_/A VGND VGND VPWR VPWR _18427_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11731__D _11731_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18358_ _18358_/A VGND VGND VPWR VPWR _18358_/Y sky130_fd_sc_hd__inv_2
X_17309_ _17254_/X _17320_/B VGND VGND VPWR VPWR _17309_/X sky130_fd_sc_hd__or2_4
XFILLER_33_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18289_ _17713_/X _18319_/B _18287_/X VGND VGND VPWR VPWR _24203_/D sky130_fd_sc_hd__o21a_4
X_20320_ _17448_/X _22389_/B VGND VGND VPWR VPWR _20320_/X sky130_fd_sc_hd__or2_4
XFILLER_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20251_ _23436_/Q VGND VGND VPWR VPWR _22367_/B sky130_fd_sc_hd__inv_2
XFILLER_115_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20182_ _20182_/A VGND VGND VPWR VPWR _20182_/X sky130_fd_sc_hd__buf_2
XFILLER_66_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24448__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11756__A _11756_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24990_ _24984_/CLK _24990_/D HRESETn VGND VGND VPWR VPWR _24990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24111__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23941_ _25122_/CLK _23941_/D HRESETn VGND VGND VPWR VPWR _18879_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_69_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23872_ _25485_/CLK _19028_/X VGND VGND VPWR VPWR _23872_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24030__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23325__A2 _22467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22823_ _12286_/B _22820_/X _22822_/X VGND VGND VPWR VPWR _22823_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__16059__A _24709_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22533__B1 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22754_ _17756_/A _22821_/A _12249_/X _22429_/A VGND VGND VPWR VPWR _22754_/X sky130_fd_sc_hd__o22a_4
X_21705_ _17244_/Y _21303_/X _25358_/Q _23100_/A VGND VGND VPWR VPWR _21706_/B sky130_fd_sc_hd__a2bb2o_4
X_25473_ _25141_/CLK _25473_/D HRESETn VGND VGND VPWR VPWR _12063_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25236__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22685_ _12238_/X _22714_/A _17755_/Y _22684_/X VGND VGND VPWR VPWR _22685_/X sky130_fd_sc_hd__o22a_4
XFILLER_9_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17960__B1 _14620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24424_ _24457_/CLK _24424_/D HRESETn VGND VGND VPWR VPWR _24424_/Q sky130_fd_sc_hd__dfrtp_4
X_21636_ _21498_/A VGND VGND VPWR VPWR _21636_/X sky130_fd_sc_hd__buf_2
X_24355_ _24355_/CLK _17286_/X HRESETn VGND VGND VPWR VPWR _24355_/Q sky130_fd_sc_hd__dfrtp_4
X_21567_ _21560_/X _21563_/X _21564_/X _21566_/X VGND VGND VPWR VPWR _21567_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17712__B1 _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23306_ _23306_/A _23305_/X VGND VGND VPWR VPWR _23313_/C sky130_fd_sc_hd__and2_4
X_20518_ _14279_/A _20504_/C _20516_/Y _20517_/X VGND VGND VPWR VPWR _20519_/B sky130_fd_sc_hd__a211o_4
X_21498_ _21498_/A _21497_/X VGND VGND VPWR VPWR _21498_/X sky130_fd_sc_hd__or2_4
XFILLER_14_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24286_ _24285_/CLK _17677_/X HRESETn VGND VGND VPWR VPWR _24286_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22524__A _22524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18268__A1 _13795_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20449_ _14541_/A _20448_/Y VGND VGND VPWR VPWR _20449_/Y sky130_fd_sc_hd__nor2_4
XFILLER_118_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23312__A2_N _23309_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19465__B1 _19420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23237_ _24461_/Q _22654_/X _23172_/X VGND VGND VPWR VPWR _23237_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24871__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18428__A1_N _21322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23168_ _24528_/Q _22922_/X _22923_/X _23167_/X VGND VGND VPWR VPWR _23169_/C sky130_fd_sc_hd__a211o_4
XFILLER_79_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24800__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22119_ _13784_/C _22083_/X _22087_/X _22093_/X _22118_/X VGND VGND VPWR VPWR _22149_/B
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__23013__A1 _12252_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19217__B1 _19149_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15990_ _24734_/Q VGND VGND VPWR VPWR _15990_/Y sky130_fd_sc_hd__inv_2
X_23099_ _23143_/A _23099_/B VGND VGND VPWR VPWR _23114_/B sky130_fd_sc_hd__and2_4
XANTENNA__24118__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14941_ _24418_/Q VGND VGND VPWR VPWR _14941_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23355__A _23342_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17660_ _17660_/A VGND VGND VPWR VPWR _17660_/Y sky130_fd_sc_hd__inv_2
X_14872_ _14798_/B _14872_/B VGND VGND VPWR VPWR _14872_/Y sky130_fd_sc_hd__nor2_4
XFILLER_85_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16611_ _16611_/A VGND VGND VPWR VPWR _16611_/Y sky130_fd_sc_hd__inv_2
X_13823_ _22726_/A _13822_/X _11800_/X _13822_/X VGND VGND VPWR VPWR _25257_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17591_ _17585_/A _17585_/B _17586_/B _17590_/X VGND VGND VPWR VPWR _17591_/X sky130_fd_sc_hd__a211o_4
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21327__A1 _24535_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16542_ _15709_/A VGND VGND VPWR VPWR _16795_/A sky130_fd_sc_hd__buf_2
X_19330_ _19329_/Y _19325_/X _19307_/X _19311_/Y VGND VGND VPWR VPWR _23765_/D sky130_fd_sc_hd__a2bb2o_4
X_13754_ _13754_/A VGND VGND VPWR VPWR _14697_/A sky130_fd_sc_hd__inv_2
XANTENNA__16203__B1 _11764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12705_ _12595_/Y _12704_/X VGND VGND VPWR VPWR _12706_/B sky130_fd_sc_hd__or2_4
X_19261_ _21225_/B _19256_/X _18919_/X _19256_/A VGND VGND VPWR VPWR _19261_/X sky130_fd_sc_hd__a2bb2o_4
X_16473_ _24560_/Q VGND VGND VPWR VPWR _16473_/Y sky130_fd_sc_hd__inv_2
X_13685_ _13685_/A _13685_/B VGND VGND VPWR VPWR _13685_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18184__A _18184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18212_ _18180_/A _23861_/Q VGND VGND VPWR VPWR _18213_/C sky130_fd_sc_hd__or2_4
X_15424_ _15092_/Y _15316_/X _15318_/A _15421_/Y VGND VGND VPWR VPWR _15425_/A sky130_fd_sc_hd__a211o_4
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12636_ _12636_/A _12636_/B VGND VGND VPWR VPWR _12637_/C sky130_fd_sc_hd__or2_4
X_19192_ _19190_/Y _19188_/X _19191_/X _19188_/X VGND VGND VPWR VPWR _19192_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21322__B _22298_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_156_0_HCLK clkbuf_7_78_0_HCLK/X VGND VGND VPWR VPWR _24275_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18143_ _18175_/A _18980_/A VGND VGND VPWR VPWR _18144_/C sky130_fd_sc_hd__or2_4
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ _24984_/Q _15355_/B VGND VGND VPWR VPWR _15357_/B sky130_fd_sc_hd__or2_4
XFILLER_8_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12567_ _12567_/A VGND VGND VPWR VPWR _12567_/Y sky130_fd_sc_hd__inv_2
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24959__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14306_ _14305_/Y VGND VGND VPWR VPWR _14306_/X sky130_fd_sc_hd__buf_2
XFILLER_106_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18074_ _17990_/A VGND VGND VPWR VPWR _18175_/A sky130_fd_sc_hd__buf_2
X_15286_ _15285_/X VGND VGND VPWR VPWR _15315_/A sky130_fd_sc_hd__inv_2
X_12498_ _12280_/Y _12509_/B VGND VGND VPWR VPWR _12499_/B sky130_fd_sc_hd__or2_4
X_17025_ _17005_/Y _17025_/B VGND VGND VPWR VPWR _17060_/A sky130_fd_sc_hd__or2_4
X_14237_ _14235_/Y _14236_/X _13803_/X _14236_/X VGND VGND VPWR VPWR _14237_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23252__B2 _22280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12543__A2 _12542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14168_ _14111_/X _14167_/Y _14446_/A _14111_/X VGND VGND VPWR VPWR _25200_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16893__A1_N _22183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24541__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13119_ _13119_/A _13119_/B _13119_/C _13119_/D VGND VGND VPWR VPWR _13120_/D sky130_fd_sc_hd__or4_4
XFILLER_86_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19743__A _19729_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14099_ _14099_/A _14098_/X _14099_/C VGND VGND VPWR VPWR _14100_/B sky130_fd_sc_hd__or3_4
X_18976_ _18976_/A VGND VGND VPWR VPWR _18976_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17927_ _13541_/B _17914_/Y _17923_/X VGND VGND VPWR VPWR _24237_/D sky130_fd_sc_hd__o21a_4
X_17858_ _17858_/A VGND VGND VPWR VPWR _24255_/D sky130_fd_sc_hd__inv_2
XFILLER_66_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16809_ _16809_/A VGND VGND VPWR VPWR _16809_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21318__A1 _24434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17789_ _17761_/X _17771_/B _17762_/A VGND VGND VPWR VPWR _17790_/C sky130_fd_sc_hd__o21a_4
XFILLER_130_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19528_ _19528_/A VGND VGND VPWR VPWR _19528_/X sky130_fd_sc_hd__buf_2
XANTENNA__16201__A1_N _16199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12200__A _22853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_52_0_HCLK clkbuf_7_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19459_ _19446_/Y VGND VGND VPWR VPWR _19459_/X sky130_fd_sc_hd__buf_2
XANTENNA__15511__A _15490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22470_ _23034_/A VGND VGND VPWR VPWR _22470_/X sky130_fd_sc_hd__buf_2
X_21421_ _22287_/A _21420_/X VGND VGND VPWR VPWR _21421_/Y sky130_fd_sc_hd__nand2_4
XFILLER_72_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19695__B1 _19599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13031__A _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21352_ _21352_/A VGND VGND VPWR VPWR _21352_/X sky130_fd_sc_hd__buf_2
X_24140_ _24136_/CLK _24140_/D HRESETn VGND VGND VPWR VPWR _18719_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_11_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20303_ _20303_/A VGND VGND VPWR VPWR _22028_/B sky130_fd_sc_hd__inv_2
XANTENNA__24629__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21283_ _22138_/A VGND VGND VPWR VPWR _21284_/A sky130_fd_sc_hd__buf_2
X_24071_ _24070_/CLK _24071_/D HRESETn VGND VGND VPWR VPWR _20505_/C sky130_fd_sc_hd__dfrtp_4
X_20234_ _20230_/Y _20233_/X _18247_/X _20233_/X VGND VGND VPWR VPWR _20234_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12534__A2 _12533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23022_ _22819_/X _23013_/Y _23017_/Y _23021_/X VGND VGND VPWR VPWR _23030_/C sky130_fd_sc_hd__a211o_4
XANTENNA__19998__B2 _19991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24282__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20165_ _20165_/A VGND VGND VPWR VPWR _20165_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24211__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16681__B1 _16325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20096_ _20096_/A VGND VGND VPWR VPWR _20096_/X sky130_fd_sc_hd__buf_2
X_24973_ _24977_/CLK _24973_/D HRESETn VGND VGND VPWR VPWR _24973_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21557__B2 _16723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22754__B1 _12249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17498__A2_N _24294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23924_ _25098_/CLK _23924_/D HRESETn VGND VGND VPWR VPWR _22161_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25488__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23855_ _23854_/CLK _19078_/X VGND VGND VPWR VPWR _13369_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16984__A1 _24712_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25417__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22806_ _22792_/Y _23002_/A _22806_/C _22806_/D VGND VGND VPWR VPWR _22806_/X sky130_fd_sc_hd__or4_4
XFILLER_38_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23786_ _24396_/CLK _23786_/D VGND VGND VPWR VPWR _23786_/Q sky130_fd_sc_hd__dfxtp_4
X_20998_ _23964_/Q VGND VGND VPWR VPWR _21000_/B sky130_fd_sc_hd__inv_2
XANTENNA__25118__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25525_ _25526_/CLK _11789_/X HRESETn VGND VGND VPWR VPWR _25525_/Q sky130_fd_sc_hd__dfrtp_4
X_22737_ _24787_/Q _22587_/B VGND VGND VPWR VPWR _22737_/X sky130_fd_sc_hd__or2_4
XFILLER_0_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25070__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13470_ _13533_/A _13533_/B _15652_/D _12059_/X VGND VGND VPWR VPWR _13471_/A sky130_fd_sc_hd__or4_4
X_25456_ _24102_/CLK _12124_/X HRESETn VGND VGND VPWR VPWR _25456_/Q sky130_fd_sc_hd__dfrtp_4
X_22668_ _22441_/X _22665_/X _22444_/X _22667_/X VGND VGND VPWR VPWR _22669_/A sky130_fd_sc_hd__o22a_4
Xclkbuf_8_229_0_HCLK clkbuf_8_229_0_HCLK/A VGND VGND VPWR VPWR _24821_/CLK sky130_fd_sc_hd__clkbuf_1
X_12421_ _12277_/B _12415_/X _12402_/X _12417_/Y VGND VGND VPWR VPWR _12422_/A sky130_fd_sc_hd__a211o_4
X_24407_ _24407_/CLK _16845_/X HRESETn VGND VGND VPWR VPWR _14890_/A sky130_fd_sc_hd__dfrtp_4
X_21619_ _21631_/A _21619_/B _21619_/C VGND VGND VPWR VPWR _21619_/X sky130_fd_sc_hd__and3_4
XFILLER_107_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25387_ _24804_/CLK _25387_/D HRESETn VGND VGND VPWR VPWR _21005_/A sky130_fd_sc_hd__dfrtp_4
X_22599_ _21105_/A _22597_/X _22103_/X _22598_/X VGND VGND VPWR VPWR _22600_/B sky130_fd_sc_hd__o22a_4
XFILLER_12_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21870__A1_N _22425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15140_ _15139_/Y _24582_/Q _15139_/Y _24582_/Q VGND VGND VPWR VPWR _15140_/X sky130_fd_sc_hd__a2bb2o_4
X_12352_ _25335_/Q VGND VGND VPWR VPWR _12352_/Y sky130_fd_sc_hd__inv_2
X_24338_ _24177_/CLK _17357_/Y HRESETn VGND VGND VPWR VPWR _17174_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_103_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11769__A1_N _11766_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22254__A _21454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15071_ _15071_/A _15070_/X VGND VGND VPWR VPWR _15072_/B sky130_fd_sc_hd__or2_4
XANTENNA__23234__A1 _24530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12283_ _12209_/Y _12269_/Y _12278_/X _12283_/D VGND VGND VPWR VPWR _12283_/X sky130_fd_sc_hd__or4_4
XANTENNA__23069__B _23069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24269_ _24692_/CLK _17800_/Y HRESETn VGND VGND VPWR VPWR _24269_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14022_ _14003_/C VGND VGND VPWR VPWR _14022_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13722__A1 _13686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22588__A3 _22127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22993__B1 _22798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18830_ _16539_/Y _18614_/X _16539_/Y _18614_/X VGND VGND VPWR VPWR _18830_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16672__B1 _16403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23085__A _23085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15973_ _15966_/X _15969_/X _11812_/X _24747_/Q _15967_/X VGND VGND VPWR VPWR _24747_/D
+ sky130_fd_sc_hd__a32o_4
X_18761_ _24130_/Q _18760_/Y VGND VGND VPWR VPWR _18761_/X sky130_fd_sc_hd__or2_4
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14924_ _14924_/A _14917_/X _14920_/X _14923_/X VGND VGND VPWR VPWR _14940_/C sky130_fd_sc_hd__or4_4
X_17712_ _21467_/A _17711_/X _21467_/A _17711_/X VGND VGND VPWR VPWR _17733_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18692_ _18692_/A _18692_/B _18692_/C _18691_/X VGND VGND VPWR VPWR _18693_/B sky130_fd_sc_hd__or4_4
XFILLER_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16424__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23934__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14855_ _14814_/C _14799_/X _14814_/C _14799_/X VGND VGND VPWR VPWR _14855_/X sky130_fd_sc_hd__a2bb2o_4
X_17643_ _17525_/Y _17639_/X VGND VGND VPWR VPWR _17643_/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15778__A2 _15655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16975__B2 _17038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13806_ _25259_/Q VGND VGND VPWR VPWR _21366_/A sky130_fd_sc_hd__inv_2
X_17574_ _24289_/Q VGND VGND VPWR VPWR _17574_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14786_ _17980_/A VGND VGND VPWR VPWR _18177_/A sky130_fd_sc_hd__buf_2
X_11998_ _11992_/B VGND VGND VPWR VPWR _11998_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22429__A _22429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16525_ _15623_/A VGND VGND VPWR VPWR _16525_/X sky130_fd_sc_hd__buf_2
X_19313_ _19017_/X VGND VGND VPWR VPWR _19313_/X sky130_fd_sc_hd__buf_2
XANTENNA__21333__A _21333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13737_ _13757_/B VGND VGND VPWR VPWR _13748_/A sky130_fd_sc_hd__buf_2
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_39_0_HCLK clkbuf_5_19_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_79_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16456_ _18496_/A _16455_/X _16366_/X _16455_/X VGND VGND VPWR VPWR _24566_/D sky130_fd_sc_hd__a2bb2o_4
X_19244_ _19256_/A VGND VGND VPWR VPWR _19244_/X sky130_fd_sc_hd__buf_2
X_13668_ _24060_/Q _13667_/X VGND VGND VPWR VPWR _13668_/X sky130_fd_sc_hd__or2_4
X_15407_ _15285_/X VGND VGND VPWR VPWR _15407_/X sky130_fd_sc_hd__buf_2
XFILLER_73_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12619_ _12611_/X _12618_/X VGND VGND VPWR VPWR _12619_/X sky130_fd_sc_hd__or2_4
X_19175_ _19175_/A VGND VGND VPWR VPWR _19175_/Y sky130_fd_sc_hd__inv_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16387_ _15090_/Y _16382_/X _16386_/X _16382_/X VGND VGND VPWR VPWR _24594_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19677__B1 _19553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13599_ _13598_/X VGND VGND VPWR VPWR _14659_/A sky130_fd_sc_hd__buf_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12359__A2_N _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24793__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18126_ _18056_/A _19208_/A VGND VGND VPWR VPWR _18126_/X sky130_fd_sc_hd__or2_4
XFILLER_8_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15338_ _15338_/A _15338_/B VGND VGND VPWR VPWR _15338_/X sky130_fd_sc_hd__or2_4
XANTENNA__24722__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18057_ _18057_/A _18057_/B _18056_/X VGND VGND VPWR VPWR _18057_/X sky130_fd_sc_hd__and3_4
XANTENNA__17258__A _17236_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15269_ _15250_/A _15267_/X _15268_/Y VGND VGND VPWR VPWR _15269_/X sky130_fd_sc_hd__o21a_4
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19429__B1 _19404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17008_ _16009_/Y _17026_/A _24723_/Q _17007_/Y VGND VGND VPWR VPWR _17008_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18959_ _18959_/A VGND VGND VPWR VPWR _18959_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21539__A1 _21275_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21970_ _21264_/X _21968_/X _21969_/X _18259_/Y _21636_/X VGND VGND VPWR VPWR _21970_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_6_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14410__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16415__B1 _16325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20921_ _20920_/X VGND VGND VPWR VPWR _24052_/D sky130_fd_sc_hd__inv_2
XANTENNA__25510__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18817__A _18682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13026__A _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23640_ _23649_/CLK _19695_/X VGND VGND VPWR VPWR _23640_/Q sky130_fd_sc_hd__dfxtp_4
X_20852_ _20846_/Y _20852_/B _20851_/Y VGND VGND VPWR VPWR _20852_/X sky130_fd_sc_hd__and3_4
XPHY_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17529__A1_N _11860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23571_ _23580_/CLK _23571_/D VGND VGND VPWR VPWR _23571_/Q sky130_fd_sc_hd__dfxtp_4
X_20783_ _24021_/Q _20783_/B VGND VGND VPWR VPWR _20783_/Y sky130_fd_sc_hd__nor2_4
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21711__B2 _17416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25310_ _25309_/CLK _13480_/X HRESETn VGND VGND VPWR VPWR _25310_/Q sky130_fd_sc_hd__dfrtp_4
X_22522_ _24577_/Q _22522_/B VGND VGND VPWR VPWR _22530_/B sky130_fd_sc_hd__or2_4
XFILLER_74_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25241_ _24148_/CLK _25241_/D HRESETn VGND VGND VPWR VPWR _13853_/A sky130_fd_sc_hd__dfrtp_4
X_22453_ _22613_/B _22451_/X _13813_/B _22452_/X VGND VGND VPWR VPWR _22453_/X sky130_fd_sc_hd__o22a_4
X_21404_ _21162_/X _21388_/X _21403_/X VGND VGND VPWR VPWR _21404_/X sky130_fd_sc_hd__and3_4
X_25172_ _25172_/CLK _25172_/D HRESETn VGND VGND VPWR VPWR _25172_/Q sky130_fd_sc_hd__dfrtp_4
X_22384_ _22384_/A VGND VGND VPWR VPWR _22384_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24463__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_59_0_HCLK clkbuf_8_59_0_HCLK/A VGND VGND VPWR VPWR _25279_/CLK sky130_fd_sc_hd__clkbuf_1
X_24123_ _24136_/CLK _18794_/Y HRESETn VGND VGND VPWR VPWR _24123_/Q sky130_fd_sc_hd__dfrtp_4
X_21335_ _21335_/A VGND VGND VPWR VPWR _21336_/A sky130_fd_sc_hd__buf_2
XFILLER_108_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24054_ _24447_/CLK _20928_/X HRESETn VGND VGND VPWR VPWR _24054_/Q sky130_fd_sc_hd__dfrtp_4
X_21266_ _22575_/A _21265_/X _13848_/Y _22575_/A VGND VGND VPWR VPWR _21266_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21778__B2 _22390_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23005_ _24556_/Q _22810_/X _23005_/C VGND VGND VPWR VPWR _23005_/X sky130_fd_sc_hd__and3_4
X_20217_ _20211_/Y VGND VGND VPWR VPWR _20217_/X sky130_fd_sc_hd__buf_2
X_21197_ _21162_/X _21180_/X _21196_/X VGND VGND VPWR VPWR _21197_/X sky130_fd_sc_hd__and3_4
XFILLER_133_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16654__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20148_ _20148_/A VGND VGND VPWR VPWR _20161_/A sky130_fd_sc_hd__inv_2
X_12970_ _12976_/A _12979_/B VGND VGND VPWR VPWR _12970_/X sky130_fd_sc_hd__or2_4
X_20079_ _20079_/A VGND VGND VPWR VPWR _20079_/X sky130_fd_sc_hd__buf_2
X_24956_ _24957_/CLK _15447_/X HRESETn VGND VGND VPWR VPWR _13920_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11921_ _11916_/A _11919_/Y _11920_/Y VGND VGND VPWR VPWR _25498_/D sky130_fd_sc_hd__o21a_4
X_23907_ _23905_/CLK _23907_/D VGND VGND VPWR VPWR _18927_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_85_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25251__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24887_ _24035_/CLK _24887_/D HRESETn VGND VGND VPWR VPWR _24887_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_72_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14640_ _18202_/A VGND VGND VPWR VPWR _18006_/A sky130_fd_sc_hd__buf_2
XFILLER_122_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11852_ _18254_/A VGND VGND VPWR VPWR _16359_/A sky130_fd_sc_hd__buf_2
X_23838_ _25488_/CLK _19123_/X VGND VGND VPWR VPWR _13402_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14571_ _14571_/A VGND VGND VPWR VPWR _14571_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17350__B _17350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11783_ _25526_/Q VGND VGND VPWR VPWR _11783_/Y sky130_fd_sc_hd__inv_2
X_23769_ _25503_/CLK _19321_/X VGND VGND VPWR VPWR _18066_/B sky130_fd_sc_hd__dfxtp_4
X_16310_ _22971_/A VGND VGND VPWR VPWR _16310_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21702__B2 _21533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13522_ _13522_/A _25167_/Q _12027_/D _13522_/D VGND VGND VPWR VPWR _13522_/X sky130_fd_sc_hd__and4_4
X_25508_ _25508_/CLK _11863_/X HRESETn VGND VGND VPWR VPWR _11860_/A sky130_fd_sc_hd__dfrtp_4
X_17290_ _17289_/X VGND VGND VPWR VPWR _24354_/D sky130_fd_sc_hd__inv_2
XFILLER_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16241_ _16225_/A VGND VGND VPWR VPWR _16241_/X sky130_fd_sc_hd__buf_2
X_13453_ _13453_/A _13451_/X _13453_/C VGND VGND VPWR VPWR _13453_/X sky130_fd_sc_hd__and3_4
X_25439_ _24759_/CLK _25439_/D HRESETn VGND VGND VPWR VPWR _12213_/A sky130_fd_sc_hd__dfrtp_4
X_12404_ _12404_/A VGND VGND VPWR VPWR _25448_/D sky130_fd_sc_hd__inv_2
X_16172_ _14769_/X _16172_/B VGND VGND VPWR VPWR _16175_/C sky130_fd_sc_hd__and2_4
X_13384_ _13316_/A _23647_/Q VGND VGND VPWR VPWR _13386_/B sky130_fd_sc_hd__or2_4
X_15123_ _24968_/Q VGND VGND VPWR VPWR _15390_/A sky130_fd_sc_hd__inv_2
XFILLER_5_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12335_ _25324_/Q _24809_/Q _13107_/A _12334_/Y VGND VGND VPWR VPWR _12335_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24133__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15054_ _15054_/A _15049_/X _15054_/C _15054_/D VGND VGND VPWR VPWR _15054_/X sky130_fd_sc_hd__or4_4
X_19931_ _19943_/A VGND VGND VPWR VPWR _19931_/X sky130_fd_sc_hd__buf_2
X_12266_ _12266_/A VGND VGND VPWR VPWR _12266_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22712__A _22266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14005_ _14042_/D VGND VGND VPWR VPWR _14005_/Y sky130_fd_sc_hd__inv_2
X_19862_ _19861_/Y _19859_/X _19797_/X _19859_/X VGND VGND VPWR VPWR _23582_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22430__A2 _22407_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12197_ _12196_/Y _24735_/Q _12196_/Y _24735_/Q VGND VGND VPWR VPWR _12198_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18634__B2 _18682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18813_ _18639_/Y _18783_/X VGND VGND VPWR VPWR _18820_/B sky130_fd_sc_hd__or2_4
X_19793_ _19793_/A VGND VGND VPWR VPWR _19793_/X sky130_fd_sc_hd__buf_2
XANTENNA__25339__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18744_ _18768_/A _18765_/A _18765_/B VGND VGND VPWR VPWR _18756_/B sky130_fd_sc_hd__or3_4
X_15956_ _12193_/Y _15954_/X _15955_/X _15954_/X VGND VGND VPWR VPWR _15956_/X sky130_fd_sc_hd__a2bb2o_4
X_14907_ _24995_/Q VGND VGND VPWR VPWR _15061_/D sky130_fd_sc_hd__inv_2
XFILLER_64_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15887_ _15857_/A VGND VGND VPWR VPWR _15887_/X sky130_fd_sc_hd__buf_2
X_18675_ _18675_/A VGND VGND VPWR VPWR _18675_/X sky130_fd_sc_hd__buf_2
X_17626_ _17568_/X _17626_/B VGND VGND VPWR VPWR _17626_/X sky130_fd_sc_hd__or2_4
XFILLER_40_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14838_ _25039_/Q _14816_/X _25039_/Q _14816_/X VGND VGND VPWR VPWR _14838_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14769_ _13588_/X VGND VGND VPWR VPWR _14769_/X sky130_fd_sc_hd__buf_2
X_17557_ _24701_/Q VGND VGND VPWR VPWR _17557_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13631__B1 _17928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24974__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16508_ _16508_/A VGND VGND VPWR VPWR _16508_/Y sky130_fd_sc_hd__inv_2
X_17488_ _13174_/X _17486_/X _13162_/X _17487_/Y VGND VGND VPWR VPWR _17488_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24903__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19227_ _19221_/Y VGND VGND VPWR VPWR _19227_/X sky130_fd_sc_hd__buf_2
XANTENNA__15996__A _15995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16439_ _24570_/Q VGND VGND VPWR VPWR _16439_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_212_0_HCLK clkbuf_8_213_0_HCLK/A VGND VGND VPWR VPWR _24596_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19158_ _19157_/Y _19154_/X _19133_/X _19154_/X VGND VGND VPWR VPWR _23827_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21510__B _21407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18109_ _14646_/X _18109_/B _18108_/X VGND VGND VPWR VPWR _18109_/X sky130_fd_sc_hd__and3_4
XFILLER_117_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19089_ _19088_/Y _19086_/X _16867_/X _19086_/X VGND VGND VPWR VPWR _19089_/X sky130_fd_sc_hd__a2bb2o_4
X_21120_ _20968_/A _14192_/X _14472_/Y _21355_/A VGND VGND VPWR VPWR _21125_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22957__B1 _11780_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21051_ _21051_/A _21026_/B VGND VGND VPWR VPWR _21059_/B sky130_fd_sc_hd__or2_4
XANTENNA__18827__A1_N _16469_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16620__A _16620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20002_ _20014_/A VGND VGND VPWR VPWR _20002_/X sky130_fd_sc_hd__buf_2
XANTENNA__12236__A2_N _24747_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22709__B1 _21103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11764__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24810_ _24842_/CLK _15838_/X HRESETn VGND VGND VPWR VPWR _24810_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22185__A1 _25513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25009__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12122__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24741_ _24792_/CLK _15981_/X HRESETn VGND VGND VPWR VPWR _22267_/A sky130_fd_sc_hd__dfrtp_4
X_21953_ _21953_/A _21362_/X VGND VGND VPWR VPWR _21953_/X sky130_fd_sc_hd__or2_4
XFILLER_41_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20904_ _20904_/A VGND VGND VPWR VPWR _20904_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24672_ _24606_/CLK _24672_/D HRESETn VGND VGND VPWR VPWR _24672_/Q sky130_fd_sc_hd__dfrtp_4
X_21884_ _21879_/X _21883_/X _14712_/A VGND VGND VPWR VPWR _21884_/X sky130_fd_sc_hd__o21a_4
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _23623_/CLK _19744_/X VGND VGND VPWR VPWR _13392_/B sky130_fd_sc_hd__dfxtp_4
X_20835_ _20834_/X VGND VGND VPWR VPWR _20835_/Y sky130_fd_sc_hd__inv_2
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16067__A _15995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23283__A1_N _17235_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_22_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23554_ _23545_/CLK _19937_/X VGND VGND VPWR VPWR _19935_/A sky130_fd_sc_hd__dfxtp_4
X_20766_ _13120_/B VGND VGND VPWR VPWR _20767_/A sky130_fd_sc_hd__inv_2
XFILLER_11_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24644__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22505_ _22505_/A VGND VGND VPWR VPWR _22505_/X sky130_fd_sc_hd__buf_2
XANTENNA__19378__A _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23485_ _23453_/CLK _23485_/D VGND VGND VPWR VPWR _23485_/Q sky130_fd_sc_hd__dfxtp_4
X_20697_ _20697_/A VGND VGND VPWR VPWR _20697_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25224_ _23967_/CLK _14077_/X HRESETn VGND VGND VPWR VPWR _13997_/A sky130_fd_sc_hd__dfrtp_4
X_22436_ _17846_/X _22425_/X _25363_/Q _22435_/X VGND VGND VPWR VPWR _22436_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25155_ _24109_/CLK _14332_/X HRESETn VGND VGND VPWR VPWR _25155_/Q sky130_fd_sc_hd__dfrtp_4
X_22367_ _22070_/X _22367_/B VGND VGND VPWR VPWR _22367_/X sky130_fd_sc_hd__or2_4
XFILLER_108_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12120_ _12118_/Y _12114_/X _11858_/X _12119_/X VGND VGND VPWR VPWR _25458_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24106_ _25205_/CLK _24106_/D HRESETn VGND VGND VPWR VPWR _24106_/Q sky130_fd_sc_hd__dfstp_4
X_21318_ _24434_/Q _21293_/X _22885_/A VGND VGND VPWR VPWR _21318_/X sky130_fd_sc_hd__o21a_4
XANTENNA__20924__A1_N _20909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25086_ _24322_/CLK _25086_/D HRESETn VGND VGND VPWR VPWR _25086_/Q sky130_fd_sc_hd__dfrtp_4
X_22298_ _15105_/A _22298_/B VGND VGND VPWR VPWR _22301_/B sky130_fd_sc_hd__or2_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12051_ _11716_/A VGND VGND VPWR VPWR _15700_/C sky130_fd_sc_hd__buf_2
X_24037_ _24581_/CLK _24037_/D HRESETn VGND VGND VPWR VPWR _20851_/A sky130_fd_sc_hd__dfrtp_4
X_21249_ _21249_/A _20186_/Y VGND VGND VPWR VPWR _21250_/C sky130_fd_sc_hd__or2_4
XANTENNA__19813__B1 _19740_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16530__A _21837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23066__C _23066_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25432__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15810_ _12308_/Y _15809_/X _11778_/X _15809_/X VGND VGND VPWR VPWR _24828_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16790_ _24434_/Q VGND VGND VPWR VPWR _16790_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15741_ _15728_/X _15713_/X _15739_/X _24858_/Q _15740_/X VGND VGND VPWR VPWR _24858_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23363__A _21006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12953_ _12955_/B VGND VGND VPWR VPWR _12953_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20187__B1 _20123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24939_ _24148_/CLK _24939_/D HRESETn VGND VGND VPWR VPWR _14876_/A sky130_fd_sc_hd__dfstp_4
XFILLER_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_104_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_104_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11904_ _11904_/A VGND VGND VPWR VPWR _11904_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17361__A _17350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15672_ _22520_/A VGND VGND VPWR VPWR _22884_/B sky130_fd_sc_hd__buf_2
X_18460_ _18460_/A _18460_/B VGND VGND VPWR VPWR _18479_/C sky130_fd_sc_hd__or2_4
XANTENNA__23082__B _23082_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12884_ _12884_/A _12879_/B _12883_/X VGND VGND VPWR VPWR _12884_/X sky130_fd_sc_hd__or3_4
X_14623_ _14614_/X _14630_/B _14622_/Y VGND VGND VPWR VPWR _14623_/X sky130_fd_sc_hd__a21o_4
X_17411_ _24068_/Q _13967_/Y _21000_/A _13886_/X VGND VGND VPWR VPWR _17411_/X sky130_fd_sc_hd__o22a_4
X_11835_ _25513_/Q VGND VGND VPWR VPWR _11835_/Y sky130_fd_sc_hd__inv_2
X_18391_ _16240_/Y _24156_/Q _16240_/Y _24156_/Q VGND VGND VPWR VPWR _18391_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17249_/Y _17336_/X _17289_/A _17338_/Y VGND VGND VPWR VPWR _17342_/X sky130_fd_sc_hd__a211o_4
XFILLER_109_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _25085_/Q VGND VGND VPWR VPWR _14554_/Y sky130_fd_sc_hd__inv_2
X_11766_ _25531_/Q VGND VGND VPWR VPWR _11766_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21151__A2 _15852_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22707__A _23097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24385__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _25299_/Q VGND VGND VPWR VPWR _13505_/Y sky130_fd_sc_hd__inv_2
X_17273_ _17273_/A VGND VGND VPWR VPWR _24358_/D sky130_fd_sc_hd__inv_2
XFILLER_70_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _25104_/Q VGND VGND VPWR VPWR _21708_/A sky130_fd_sc_hd__inv_2
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11697_ _24226_/Q VGND VGND VPWR VPWR _11697_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24314__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16224_ _16192_/A VGND VGND VPWR VPWR _16225_/A sky130_fd_sc_hd__buf_2
X_19012_ _23876_/Q VGND VGND VPWR VPWR _19012_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16615__A1_N _16613_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13436_ _13303_/A _13436_/B VGND VGND VPWR VPWR _13436_/X sky130_fd_sc_hd__or2_4
XANTENNA__21330__B _21350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22100__B2 _22111_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11927__B1 RsRx_S1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16155_ _16154_/Y _16152_/X _16064_/X _16152_/X VGND VGND VPWR VPWR _16155_/X sky130_fd_sc_hd__a2bb2o_4
X_13367_ _13200_/X _13351_/X _13366_/X _25317_/Q _11965_/X VGND VGND VPWR VPWR _13367_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__18855__B2 _18789_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15106_ _24970_/Q _15105_/A _15392_/A _15105_/Y VGND VGND VPWR VPWR _15106_/X sky130_fd_sc_hd__o22a_4
X_12318_ _24815_/Q VGND VGND VPWR VPWR _12318_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_42_0_HCLK clkbuf_8_43_0_HCLK/A VGND VGND VPWR VPWR _23722_/CLK sky130_fd_sc_hd__clkbuf_1
X_16086_ _16086_/A VGND VGND VPWR VPWR _16087_/A sky130_fd_sc_hd__buf_2
X_13298_ _13440_/A _23857_/Q VGND VGND VPWR VPWR _13298_/X sky130_fd_sc_hd__or2_4
XANTENNA__21984__C _21875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22442__A _23069_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15037_ _15250_/A _24440_/Q _15250_/A _24440_/Q VGND VGND VPWR VPWR _15037_/X sky130_fd_sc_hd__a2bb2o_4
X_19914_ _19913_/Y _19911_/X _19780_/X _19911_/X VGND VGND VPWR VPWR _19914_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12249_ _12248_/Y VGND VGND VPWR VPWR _12249_/X sky130_fd_sc_hd__buf_2
XFILLER_130_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23257__B _23019_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19804__B1 _18247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24942__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19845_ _19844_/X _13762_/X _19845_/C VGND VGND VPWR VPWR _19846_/A sky130_fd_sc_hd__or3_4
XFILLER_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17255__B _17249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19776_ _19793_/A VGND VGND VPWR VPWR _19776_/X sky130_fd_sc_hd__buf_2
XANTENNA__25102__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16988_ _16029_/A _16987_/A _16029_/Y _17034_/A VGND VGND VPWR VPWR _16988_/X sky130_fd_sc_hd__o22a_4
XFILLER_84_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21208__D _21207_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18727_ _18673_/Y _18736_/A VGND VGND VPWR VPWR _18728_/B sky130_fd_sc_hd__or2_4
X_15939_ _15938_/X VGND VGND VPWR VPWR _15939_/X sky130_fd_sc_hd__buf_2
XFILLER_114_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20178__B1 _20089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18658_ _18658_/A VGND VGND VPWR VPWR _18658_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23116__B1 _12749_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17609_ _17885_/B _17604_/Y _17608_/X VGND VGND VPWR VPWR _17609_/X sky130_fd_sc_hd__or3_4
XFILLER_36_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18589_ _18589_/A _18589_/B _18582_/C VGND VGND VPWR VPWR _24148_/D sky130_fd_sc_hd__and3_4
XANTENNA__12846__C _12944_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20620_ _20620_/A _20620_/B VGND VGND VPWR VPWR _20621_/B sky130_fd_sc_hd__nand2_4
XFILLER_20_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20551_ _20551_/A VGND VGND VPWR VPWR _20551_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14450__A1_N _14177_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24055__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23270_ _23095_/X _23269_/X _23141_/X _24837_/Q _23097_/X VGND VGND VPWR VPWR _23271_/B
+ sky130_fd_sc_hd__a32o_4
X_20482_ _14205_/Y _15449_/A _20480_/X _15449_/A _20481_/X VGND VGND VPWR VPWR _20483_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_118_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22221_ _23691_/Q _21995_/Y _22506_/B _22220_/X VGND VGND VPWR VPWR _22222_/A sky130_fd_sc_hd__a211o_4
XANTENNA__11759__A _25533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20102__B1 _19841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24037__CLK _24581_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22152_ _14890_/A _21312_/X _22997_/A _22151_/X VGND VGND VPWR VPWR _22153_/C sky130_fd_sc_hd__a211o_4
XFILLER_105_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21103_ _21103_/A VGND VGND VPWR VPWR _21103_/X sky130_fd_sc_hd__buf_2
X_22083_ _21260_/X _22044_/Y _22049_/X _21502_/A _22082_/X VGND VGND VPWR VPWR _22083_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_102_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21034_ _21034_/A VGND VGND VPWR VPWR _21034_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22985_ _22985_/A _23052_/B VGND VGND VPWR VPWR _22985_/X sky130_fd_sc_hd__and2_4
XANTENNA__24896__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24724_ _24715_/CLK _16023_/X HRESETn VGND VGND VPWR VPWR _24724_/Q sky130_fd_sc_hd__dfrtp_4
X_21936_ _17706_/A _21934_/X _21935_/X VGND VGND VPWR VPWR _21936_/X sky130_fd_sc_hd__and3_4
XFILLER_43_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24825__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15596__B1 _11791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24655_ _24517_/CLK _16213_/X HRESETn VGND VGND VPWR VPWR _22992_/A sky130_fd_sc_hd__dfrtp_4
X_21867_ _21085_/A VGND VGND VPWR VPWR _22644_/B sky130_fd_sc_hd__buf_2
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12743__A2_N _24783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _23478_/CLK _19798_/X VGND VGND VPWR VPWR _19796_/A sky130_fd_sc_hd__dfxtp_4
X_20818_ _20909_/A VGND VGND VPWR VPWR _20818_/X sky130_fd_sc_hd__buf_2
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24586_ _24596_/CLK _24586_/D HRESETn VGND VGND VPWR VPWR _15096_/A sky130_fd_sc_hd__dfrtp_4
X_21798_ _21794_/X _21797_/X _18299_/X VGND VGND VPWR VPWR _21799_/C sky130_fd_sc_hd__o21a_4
XANTENNA__18534__B1 _18487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23537_ _23714_/CLK _19986_/X VGND VGND VPWR VPWR _19984_/A sky130_fd_sc_hd__dfxtp_4
X_20749_ _13119_/C VGND VGND VPWR VPWR _20749_/Y sky130_fd_sc_hd__inv_2
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16525__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22881__A2 _21067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _25174_/Q VGND VGND VPWR VPWR _21548_/A sky130_fd_sc_hd__inv_2
XANTENNA__21150__B _15852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23468_ _23516_/CLK _23468_/D VGND VGND VPWR VPWR _23468_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13221_ _13212_/A VGND VGND VPWR VPWR _13270_/A sky130_fd_sc_hd__buf_2
X_25207_ _25205_/CLK _25207_/D HRESETn VGND VGND VPWR VPWR _14102_/A sky130_fd_sc_hd__dfrtp_4
X_22419_ _22419_/A VGND VGND VPWR VPWR _22419_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18837__B2 _18682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23399_ _24923_/CLK _23399_/D VGND VGND VPWR VPWR _23399_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_124_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13152_ _13248_/A VGND VGND VPWR VPWR _13180_/A sky130_fd_sc_hd__buf_2
XANTENNA__23358__A _20984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_1_0_HCLK clkbuf_8_1_0_HCLK/A VGND VGND VPWR VPWR _24396_/CLK sky130_fd_sc_hd__clkbuf_1
X_25138_ _24943_/CLK _25138_/D HRESETn VGND VGND VPWR VPWR _25138_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_29_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12103_ _12092_/Y _12102_/X _11825_/X _12102_/X VGND VGND VPWR VPWR _12103_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13083_ _12377_/Y _13082_/X VGND VGND VPWR VPWR _13084_/B sky130_fd_sc_hd__or2_4
X_17960_ _15677_/X _15684_/A _14620_/A _15918_/X VGND VGND VPWR VPWR _17960_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15520__B1 HADDR[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25069_ _25054_/CLK _25069_/D HRESETn VGND VGND VPWR VPWR _14626_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22397__A1 _11831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12034_ _12034_/A VGND VGND VPWR VPWR _12034_/X sky130_fd_sc_hd__buf_2
X_16911_ _24252_/Q VGND VGND VPWR VPWR _16911_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23929__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17891_ _17891_/A VGND VGND VPWR VPWR _17891_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19630_ _19627_/Y _19628_/X _19629_/X _19628_/X VGND VGND VPWR VPWR _19630_/X sky130_fd_sc_hd__a2bb2o_4
X_16842_ _14916_/Y _16840_/X _16604_/X _16840_/X VGND VGND VPWR VPWR _16842_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_24_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19561_ _19561_/A VGND VGND VPWR VPWR _19574_/A sky130_fd_sc_hd__inv_2
X_13985_ _25216_/Q _13985_/B VGND VGND VPWR VPWR _14003_/B sky130_fd_sc_hd__or2_4
X_16773_ _16773_/A VGND VGND VPWR VPWR _16773_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13834__B1 _11829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18512_ _18460_/A _18514_/B _18511_/Y VGND VGND VPWR VPWR _18512_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17091__A _17023_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12936_ _12936_/A _12934_/X _12935_/X VGND VGND VPWR VPWR _25368_/D sky130_fd_sc_hd__and3_4
X_15724_ _15548_/X _15713_/X _15723_/X _24868_/Q _15711_/X VGND VGND VPWR VPWR _15724_/X
+ sky130_fd_sc_hd__a32o_4
X_19492_ _17708_/Y _19492_/B _17713_/X VGND VGND VPWR VPWR _19492_/X sky130_fd_sc_hd__or3_4
XFILLER_37_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24566__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18443_ _23004_/A _18442_/Y _16214_/Y _24165_/Q VGND VGND VPWR VPWR _18444_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12867_ _12830_/Y _12864_/X _12858_/Y _12866_/X VGND VGND VPWR VPWR _12868_/A sky130_fd_sc_hd__a211o_4
X_15655_ _15655_/A VGND VGND VPWR VPWR _15655_/X sky130_fd_sc_hd__buf_2
XFILLER_61_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11818_ _11818_/A VGND VGND VPWR VPWR _11818_/X sky130_fd_sc_hd__buf_2
X_14606_ _13573_/Y _14561_/X VGND VGND VPWR VPWR _14606_/Y sky130_fd_sc_hd__nand2_4
X_15586_ _22985_/A _15581_/X _11778_/X _15581_/X VGND VGND VPWR VPWR _24901_/D sky130_fd_sc_hd__a2bb2o_4
X_18374_ _24184_/Q VGND VGND VPWR VPWR _18374_/Y sky130_fd_sc_hd__inv_2
X_12798_ _25367_/Q VGND VGND VPWR VPWR _12799_/A sky130_fd_sc_hd__inv_2
XFILLER_18_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21124__A2 _21139_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22321__A1 _22320_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12253__A1_N _12252_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _13984_/X _14536_/Y _13995_/X VGND VGND VPWR VPWR _14538_/C sky130_fd_sc_hd__o21a_4
X_17325_ _22815_/A _17324_/Y VGND VGND VPWR VPWR _17325_/X sky130_fd_sc_hd__or2_4
X_11749_ HWDATA[29] VGND VGND VPWR VPWR _11749_/X sky130_fd_sc_hd__buf_2
XANTENNA__20332__B1 _20072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ _25110_/Q VGND VGND VPWR VPWR _14468_/Y sky130_fd_sc_hd__inv_2
X_17256_ _17247_/X _17255_/X VGND VGND VPWR VPWR _17256_/X sky130_fd_sc_hd__or2_4
XANTENNA__13778__B _14406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13419_ _13246_/X _13419_/B VGND VGND VPWR VPWR _13419_/X sky130_fd_sc_hd__or2_4
X_16207_ _16207_/A VGND VGND VPWR VPWR _16207_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22085__B1 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17187_ _23073_/A _23072_/A _16302_/Y _17293_/A VGND VGND VPWR VPWR _17187_/X sky130_fd_sc_hd__o22a_4
X_14399_ _14399_/A VGND VGND VPWR VPWR _20968_/A sky130_fd_sc_hd__inv_2
XANTENNA__16839__B1 _11821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16138_ _16125_/X VGND VGND VPWR VPWR _16138_/X sky130_fd_sc_hd__buf_2
XFILLER_6_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23268__A _23245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25354__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16069_ _24706_/Q VGND VGND VPWR VPWR _16069_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12821__A1_N _12819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19828_ _19828_/A VGND VGND VPWR VPWR _19828_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21516__A _23314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19759_ _19751_/Y VGND VGND VPWR VPWR _19759_/X sky130_fd_sc_hd__buf_2
XANTENNA__16507__A1_N _16506_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22770_ _21511_/X VGND VGND VPWR VPWR _22770_/X sky130_fd_sc_hd__buf_2
X_21721_ _21714_/Y _21715_/Y _21718_/Y _21720_/Y VGND VGND VPWR VPWR _21721_/X sky130_fd_sc_hd__or4_4
XFILLER_25_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15578__B1 _11767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24236__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24440_ _24998_/CLK _16777_/X HRESETn VGND VGND VPWR VPWR _24440_/Q sky130_fd_sc_hd__dfrtp_4
X_21652_ _21460_/A _21652_/B _21652_/C VGND VGND VPWR VPWR _21652_/X sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_5_10_0_HCLK_A clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17319__A1 _17254_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22347__A _21458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21115__A2 _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20603_ _13886_/X _20602_/X _13963_/X VGND VGND VPWR VPWR _23960_/D sky130_fd_sc_hd__and3_4
X_24371_ _24364_/CLK _17137_/X HRESETn VGND VGND VPWR VPWR _24371_/Q sky130_fd_sc_hd__dfrtp_4
X_21583_ _22827_/A VGND VGND VPWR VPWR _22280_/A sky130_fd_sc_hd__buf_2
XANTENNA__12800__B2 _22623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23322_ _22792_/A _23321_/Y VGND VGND VPWR VPWR _23322_/Y sky130_fd_sc_hd__nor2_4
X_20534_ _20537_/A _20582_/B VGND VGND VPWR VPWR _20534_/X sky130_fd_sc_hd__and2_4
X_23253_ _16648_/Y _22824_/X _15565_/Y _22827_/X VGND VGND VPWR VPWR _23253_/X sky130_fd_sc_hd__o22a_4
X_20465_ _20485_/B VGND VGND VPWR VPWR _20474_/B sky130_fd_sc_hd__buf_2
X_22204_ _21388_/A _22196_/X _22203_/X VGND VGND VPWR VPWR _22204_/X sky130_fd_sc_hd__and3_4
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23184_ _24626_/Q _21519_/B VGND VGND VPWR VPWR _23184_/X sky130_fd_sc_hd__or2_4
X_20396_ _23379_/Q _20395_/Y _20976_/A _20394_/X VGND VGND VPWR VPWR _23379_/D sky130_fd_sc_hd__o22a_4
XANTENNA__25095__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22135_ _22929_/A VGND VGND VPWR VPWR _22135_/X sky130_fd_sc_hd__buf_2
XANTENNA__15502__B1 HADDR[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25024__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22066_ _22061_/X _22065_/X _14677_/X VGND VGND VPWR VPWR _22066_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_88_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22810__A _22836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21017_ _25355_/Q _21017_/B VGND VGND VPWR VPWR _21017_/X sky130_fd_sc_hd__or2_4
XFILLER_59_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23328__B1 _23172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18643__A1_N _16592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22000__B1 _21504_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13770_ _13769_/Y VGND VGND VPWR VPWR _13770_/X sky130_fd_sc_hd__buf_2
XFILLER_28_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22968_ _21416_/A VGND VGND VPWR VPWR _22968_/X sky130_fd_sc_hd__buf_2
XFILLER_83_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12721_ _12664_/A VGND VGND VPWR VPWR _12721_/X sky130_fd_sc_hd__buf_2
X_21919_ _21944_/A _19875_/Y VGND VGND VPWR VPWR _21921_/B sky130_fd_sc_hd__or2_4
XANTENNA__15569__B1 _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24707_ _24356_/CLK _16068_/X HRESETn VGND VGND VPWR VPWR _24707_/Q sky130_fd_sc_hd__dfrtp_4
X_22899_ _22899_/A _22898_/X VGND VGND VPWR VPWR _22899_/X sky130_fd_sc_hd__or2_4
X_15440_ _13957_/B _15437_/X _15432_/X _13924_/X _15438_/X VGND VGND VPWR VPWR _15440_/X
+ sky130_fd_sc_hd__a32o_4
X_12652_ _12656_/A _12656_/B VGND VGND VPWR VPWR _12652_/X sky130_fd_sc_hd__or2_4
XANTENNA__22839__C1 _22838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24638_ _24162_/CLK _16260_/X HRESETn VGND VGND VPWR VPWR _21836_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22303__B2 _21139_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ _15365_/A _15365_/B VGND VGND VPWR VPWR _15371_/Y sky130_fd_sc_hd__nand2_4
XFILLER_54_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ _12616_/B _24846_/Q _12606_/A _12582_/Y VGND VGND VPWR VPWR _12583_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20314__B1 _19995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24569_ _24465_/CLK _24569_/D HRESETn VGND VGND VPWR VPWR _15115_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14322_ _14305_/Y _14321_/X _25305_/Q _13644_/X VGND VGND VPWR VPWR _14322_/X sky130_fd_sc_hd__o22a_4
X_17110_ _17108_/A _17110_/B _17109_/Y VGND VGND VPWR VPWR _24377_/D sky130_fd_sc_hd__and3_4
XFILLER_12_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18090_ _18187_/A _19162_/A VGND VGND VPWR VPWR _18090_/X sky130_fd_sc_hd__or2_4
XFILLER_106_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23959__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13598__B _13593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17041_ _17156_/A _16985_/Y _17041_/C _17041_/D VGND VGND VPWR VPWR _17041_/X sky130_fd_sc_hd__or4_4
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ _14247_/Y _14252_/Y sda_oen_o_S5 _14247_/Y VGND VGND VPWR VPWR _25180_/D
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15741__B1 _24858_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13204_ _13440_/A _13204_/B VGND VGND VPWR VPWR _13204_/X sky130_fd_sc_hd__or2_4
X_14184_ _14184_/A VGND VGND VPWR VPWR _14184_/Y sky130_fd_sc_hd__inv_2
X_13135_ _13135_/A VGND VGND VPWR VPWR _20783_/B sky130_fd_sc_hd__buf_2
XFILLER_3_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18992_ HWDATA[6] VGND VGND VPWR VPWR _19642_/A sky130_fd_sc_hd__buf_2
X_13066_ _25337_/Q _13065_/Y VGND VGND VPWR VPWR _13066_/X sky130_fd_sc_hd__or2_4
X_17943_ _17939_/X _17942_/X _18006_/A VGND VGND VPWR VPWR _17943_/X sky130_fd_sc_hd__o21a_4
XFILLER_26_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_116_0_HCLK clkbuf_7_58_0_HCLK/X VGND VGND VPWR VPWR _24553_/CLK sky130_fd_sc_hd__clkbuf_1
X_12017_ _12015_/A _11994_/X _12016_/Y VGND VGND VPWR VPWR _12017_/X sky130_fd_sc_hd__o21a_4
XFILLER_66_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17874_ _17874_/A _17867_/B _17873_/X VGND VGND VPWR VPWR _24250_/D sky130_fd_sc_hd__and3_4
Xclkbuf_8_179_0_HCLK clkbuf_7_89_0_HCLK/X VGND VGND VPWR VPWR _24305_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23319__B1 _22786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18994__B1 _18993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19613_ _19608_/Y _19611_/X _19612_/X _19611_/X VGND VGND VPWR VPWR _23668_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24747__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16825_ _16840_/A VGND VGND VPWR VPWR _16825_/X sky130_fd_sc_hd__buf_2
XANTENNA__13807__B1 _13515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11862__A _11862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19544_ _19538_/X VGND VGND VPWR VPWR _19544_/X sky130_fd_sc_hd__buf_2
XFILLER_93_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16756_ _16755_/Y _16753_/X _16408_/X _16753_/X VGND VGND VPWR VPWR _24451_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13968_ _13968_/A VGND VGND VPWR VPWR _13969_/A sky130_fd_sc_hd__inv_2
XANTENNA__17252__C _17252_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21345__A2 _12096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22542__A1 _16597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15707_ _22123_/A VGND VGND VPWR VPWR _15708_/A sky130_fd_sc_hd__buf_2
XFILLER_46_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12919_ _12915_/X VGND VGND VPWR VPWR _12919_/Y sky130_fd_sc_hd__inv_2
X_19475_ _19475_/A VGND VGND VPWR VPWR _22020_/B sky130_fd_sc_hd__inv_2
X_13899_ _13909_/A VGND VGND VPWR VPWR _13899_/X sky130_fd_sc_hd__buf_2
X_16687_ _24479_/Q VGND VGND VPWR VPWR _16687_/Y sky130_fd_sc_hd__inv_2
X_18426_ _24146_/Q VGND VGND VPWR VPWR _18475_/C sky130_fd_sc_hd__inv_2
X_15638_ _24880_/Q VGND VGND VPWR VPWR _15638_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14232__B1 _13797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21071__A _21071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18357_ _24188_/Q _17482_/X _18356_/X VGND VGND VPWR VPWR _18358_/A sky130_fd_sc_hd__a21o_4
X_15569_ _15567_/Y _15563_/X _11754_/X _15568_/X VGND VGND VPWR VPWR _24908_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15980__B1 _15620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22845__A2 _21428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12794__B1 _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17308_ _17252_/A _17252_/B _17307_/X VGND VGND VPWR VPWR _17320_/B sky130_fd_sc_hd__or3_4
XFILLER_33_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18288_ _20000_/C _18287_/X _20000_/C _18287_/X VGND VGND VPWR VPWR _24204_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25535__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17239_ _17239_/A _17293_/A VGND VGND VPWR VPWR _17239_/X sky130_fd_sc_hd__or2_4
X_20250_ _20249_/Y _20245_/X _19771_/X _20232_/Y VGND VGND VPWR VPWR _23437_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19474__B2 _19471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20181_ _20181_/A VGND VGND VPWR VPWR _20181_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_12_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_12_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12760__A1_N _25376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14413__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_75_0_HCLK clkbuf_7_75_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_75_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21569__C1 _21568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21033__A1 _12604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23940_ _25122_/CLK _23940_/D HRESETn VGND VGND VPWR VPWR _20574_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_9_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18985__B1 _17443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24488__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23871_ _25488_/CLK _23871_/D VGND VGND VPWR VPWR _19029_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24417__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22822_ _12850_/B _21438_/X _17758_/B _22821_/X VGND VGND VPWR VPWR _22822_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14471__B1 _14470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22533__A1 _21270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22753_ _21872_/X VGND VGND VPWR VPWR _22753_/X sky130_fd_sc_hd__buf_2
XFILLER_77_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21704_ _12264_/X _22489_/A _24248_/Q _21422_/X VGND VGND VPWR VPWR _21704_/X sky130_fd_sc_hd__a2bb2o_4
X_25472_ _25309_/CLK _25472_/D HRESETn VGND VGND VPWR VPWR _12076_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23089__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22684_ _22425_/A VGND VGND VPWR VPWR _22684_/X sky130_fd_sc_hd__buf_2
XANTENNA__22077__A _22055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24423_ _24427_/CLK _24423_/D HRESETn VGND VGND VPWR VPWR _14971_/A sky130_fd_sc_hd__dfrtp_4
X_21635_ _21994_/A VGND VGND VPWR VPWR _22531_/B sky130_fd_sc_hd__buf_2
XANTENNA__15971__B1 _24749_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16075__A _16075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24354_ _24355_/CLK _24354_/D HRESETn VGND VGND VPWR VPWR _17236_/A sky130_fd_sc_hd__dfrtp_4
X_21566_ _21565_/X VGND VGND VPWR VPWR _21566_/X sky130_fd_sc_hd__buf_2
XFILLER_138_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25276__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23305_ _21863_/X _23304_/X _22466_/X _24873_/Q _21067_/A VGND VGND VPWR VPWR _23305_/X
+ sky130_fd_sc_hd__a32o_4
X_20517_ _20517_/A _20491_/A _20494_/A _20517_/D VGND VGND VPWR VPWR _20517_/X sky130_fd_sc_hd__or4_4
XFILLER_126_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24285_ _24285_/CLK _17679_/X HRESETn VGND VGND VPWR VPWR _17512_/A sky130_fd_sc_hd__dfrtp_4
X_21497_ _20333_/A _20318_/X _23381_/Q _19585_/A VGND VGND VPWR VPWR _21497_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25205__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23236_ _24595_/Q _23327_/B VGND VGND VPWR VPWR _23236_/X sky130_fd_sc_hd__or2_4
X_20448_ _25138_/Q _20446_/X _20454_/C _20447_/X VGND VGND VPWR VPWR _20448_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__23261__A2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11947__A _11947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23167_ _24560_/Q _23166_/X _23130_/X VGND VGND VPWR VPWR _23167_/X sky130_fd_sc_hd__o21a_4
X_20379_ _19536_/Y VGND VGND VPWR VPWR _20379_/X sky130_fd_sc_hd__buf_2
XFILLER_69_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22118_ _21332_/Y _22101_/X _22105_/Y _22110_/Y _22117_/X VGND VGND VPWR VPWR _22118_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23098_ _23095_/X _23096_/X _22854_/X _24832_/Q _23097_/X VGND VGND VPWR VPWR _23099_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_47_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14940_ _14940_/A _14940_/B _14940_/C _14939_/X VGND VGND VPWR VPWR _14940_/X sky130_fd_sc_hd__or4_4
X_22049_ _25247_/Q _22506_/B _13782_/X _22048_/Y VGND VGND VPWR VPWR _22049_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24840__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22772__B2 _22480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14871_ _14871_/A VGND VGND VPWR VPWR _14872_/B sky130_fd_sc_hd__buf_2
XFILLER_63_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16610_ _16608_/Y _16609_/X _16525_/X _16609_/X VGND VGND VPWR VPWR _24508_/D sky130_fd_sc_hd__a2bb2o_4
X_13822_ _13822_/A VGND VGND VPWR VPWR _13822_/X sky130_fd_sc_hd__buf_2
XFILLER_29_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17590_ _17885_/B VGND VGND VPWR VPWR _17590_/X sky130_fd_sc_hd__buf_2
XFILLER_47_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21327__A2 _22592_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13753_ _25267_/Q VGND VGND VPWR VPWR _20043_/A sky130_fd_sc_hd__buf_2
X_16541_ _16541_/A VGND VGND VPWR VPWR _16541_/Y sky130_fd_sc_hd__inv_2
X_12704_ _12704_/A _12704_/B VGND VGND VPWR VPWR _12704_/X sky130_fd_sc_hd__or2_4
X_19260_ _19260_/A VGND VGND VPWR VPWR _21225_/B sky130_fd_sc_hd__inv_2
X_13684_ _11656_/Y _13684_/B VGND VGND VPWR VPWR _13685_/B sky130_fd_sc_hd__or2_4
X_16472_ _16471_/Y _16467_/X _16386_/X _16467_/X VGND VGND VPWR VPWR _16472_/X sky130_fd_sc_hd__a2bb2o_4
X_18211_ _18211_/A _23869_/Q VGND VGND VPWR VPWR _18213_/B sky130_fd_sc_hd__or2_4
XFILLER_70_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12635_ _25417_/Q _12635_/B VGND VGND VPWR VPWR _12635_/X sky130_fd_sc_hd__or2_4
X_15423_ _15423_/A _15423_/B _15407_/X VGND VGND VPWR VPWR _24964_/D sky130_fd_sc_hd__and3_4
XFILLER_19_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19191_ _19055_/X VGND VGND VPWR VPWR _19191_/X sky130_fd_sc_hd__buf_2
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12944__C _12944_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20838__A1 _20837_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15354_ _15354_/A VGND VGND VPWR VPWR _15355_/B sky130_fd_sc_hd__inv_2
X_18142_ _17973_/X _19458_/A VGND VGND VPWR VPWR _18144_/B sky130_fd_sc_hd__or2_4
XFILLER_19_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ _12565_/Y _24854_/Q _12565_/Y _24854_/Q VGND VGND VPWR VPWR _12566_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15320__C _15310_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14305_ _13644_/X VGND VGND VPWR VPWR _14305_/Y sky130_fd_sc_hd__inv_2
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15285_ _15165_/B VGND VGND VPWR VPWR _15285_/X sky130_fd_sc_hd__buf_2
X_18073_ _18211_/A _18073_/B VGND VGND VPWR VPWR _18073_/X sky130_fd_sc_hd__or2_4
X_12497_ _12496_/X VGND VGND VPWR VPWR _12497_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14236_ _14224_/A VGND VGND VPWR VPWR _14236_/X sky130_fd_sc_hd__buf_2
X_17024_ _17023_/Y VGND VGND VPWR VPWR _17050_/A sky130_fd_sc_hd__buf_2
XFILLER_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23252__A2 _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11857__A _11856_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24999__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14167_ _14166_/X VGND VGND VPWR VPWR _14167_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14233__A _25184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13118_ _13118_/A _20790_/A VGND VGND VPWR VPWR _13118_/X sky130_fd_sc_hd__or2_4
XFILLER_98_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24928__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14098_ _14098_/A _14173_/A _25197_/Q _14098_/D VGND VGND VPWR VPWR _14098_/X sky130_fd_sc_hd__or4_4
X_18975_ _18974_/Y _18972_/X _18955_/X _18972_/X VGND VGND VPWR VPWR _23889_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13049_ _13049_/A _13047_/X _13048_/X VGND VGND VPWR VPWR _13049_/X sky130_fd_sc_hd__and3_4
X_17926_ _13541_/A _17924_/Y _17920_/C _17925_/X VGND VGND VPWR VPWR _17926_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24581__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13791__B _14255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17857_ _16898_/X _17856_/X _17790_/A _17853_/B VGND VGND VPWR VPWR _17858_/A sky130_fd_sc_hd__a211o_4
XFILLER_67_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24510__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16808_ _16806_/Y _16807_/X _15723_/X _16807_/X VGND VGND VPWR VPWR _24427_/D sky130_fd_sc_hd__a2bb2o_4
X_17788_ _17805_/A VGND VGND VPWR VPWR _17790_/A sky130_fd_sc_hd__buf_2
XFILLER_93_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15796__A3 _15714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21318__A2 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19527_ _19527_/A VGND VGND VPWR VPWR _19527_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23281__A _23281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16739_ _16739_/A VGND VGND VPWR VPWR _16739_/X sky130_fd_sc_hd__buf_2
XANTENNA__15999__A _24733_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21869__A3 _15854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19458_ _19458_/A VGND VGND VPWR VPWR _19458_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21513__B _22998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18409_ _18409_/A VGND VGND VPWR VPWR _18460_/B sky130_fd_sc_hd__inv_2
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19389_ _16786_/X VGND VGND VPWR VPWR _19389_/X sky130_fd_sc_hd__buf_2
XANTENNA__15953__B1 _15952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14408__A _11733_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21420_ _21413_/X _21414_/X _21416_/X _12562_/A _22540_/A VGND VGND VPWR VPWR _21420_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_37_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21351_ _21351_/A _21351_/B VGND VGND VPWR VPWR _21351_/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20302_ _22235_/B _20299_/X _19978_/X _20299_/X VGND VGND VPWR VPWR _23418_/D sky130_fd_sc_hd__a2bb2o_4
X_24070_ _24070_/CLK _20504_/X HRESETn VGND VGND VPWR VPWR _24070_/Q sky130_fd_sc_hd__dfstp_4
X_21282_ _21281_/X VGND VGND VPWR VPWR _22138_/A sky130_fd_sc_hd__inv_2
XFILLER_11_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11767__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23021_ _23021_/A _23021_/B _23021_/C VGND VGND VPWR VPWR _23021_/X sky130_fd_sc_hd__and3_4
X_20233_ _20232_/Y VGND VGND VPWR VPWR _20233_/X sky130_fd_sc_hd__buf_2
XANTENNA__22451__B1 _13575_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24669__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20164_ _20163_/Y _20161_/X _20099_/X _20161_/X VGND VGND VPWR VPWR _20164_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22360__A _14682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20095_ _20095_/A VGND VGND VPWR VPWR _20095_/X sky130_fd_sc_hd__buf_2
X_24972_ _24980_/CLK _24972_/D HRESETn VGND VGND VPWR VPWR _15111_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18958__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22754__B2 _22429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23923_ _23995_/CLK _23923_/D HRESETn VGND VGND VPWR VPWR _14036_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21407__C _21361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_162_0_HCLK clkbuf_7_81_0_HCLK/X VGND VGND VPWR VPWR _23394_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24251__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_5_0_HCLK clkbuf_6_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23854_ _23854_/CLK _19080_/X VGND VGND VPWR VPWR _13401_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_19_0_HCLK clkbuf_7_9_0_HCLK/X VGND VGND VPWR VPWR _24097_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22805_ _16452_/A _22802_/X _22805_/C VGND VGND VPWR VPWR _22806_/D sky130_fd_sc_hd__and3_4
XFILLER_77_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23785_ _24396_/CLK _23785_/D VGND VGND VPWR VPWR _19273_/A sky130_fd_sc_hd__dfxtp_4
X_20997_ _20996_/X VGND VGND VPWR VPWR _23964_/D sky130_fd_sc_hd__inv_2
XFILLER_26_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15702__A _15702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25524_ _25436_/CLK _25524_/D HRESETn VGND VGND VPWR VPWR _25524_/Q sky130_fd_sc_hd__dfrtp_4
X_22736_ _22736_/A _22736_/B _22736_/C VGND VGND VPWR VPWR _22736_/X sky130_fd_sc_hd__and3_4
XFILLER_77_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25457__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25455_ _24102_/CLK _25455_/D HRESETn VGND VGND VPWR VPWR _18370_/A sky130_fd_sc_hd__dfrtp_4
X_22667_ _16590_/Y _22394_/X _21573_/X _22666_/X VGND VGND VPWR VPWR _22667_/X sky130_fd_sc_hd__o22a_4
X_12420_ _12389_/A _12420_/B _12420_/C VGND VGND VPWR VPWR _12420_/X sky130_fd_sc_hd__and3_4
XFILLER_71_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24406_ _24407_/CLK _16846_/X HRESETn VGND VGND VPWR VPWR _14945_/A sky130_fd_sc_hd__dfrtp_4
X_21618_ _21618_/A _21618_/B VGND VGND VPWR VPWR _21619_/C sky130_fd_sc_hd__or2_4
X_25386_ _24780_/CLK _25386_/D HRESETn VGND VGND VPWR VPWR _12859_/A sky130_fd_sc_hd__dfrtp_4
X_22598_ _22598_/A _22598_/B VGND VGND VPWR VPWR _22598_/X sky130_fd_sc_hd__and2_4
XFILLER_138_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12351_ _12343_/X _12346_/X _12348_/X _12350_/X VGND VGND VPWR VPWR _12351_/X sky130_fd_sc_hd__or4_4
X_24337_ _24334_/CLK _24337_/D HRESETn VGND VGND VPWR VPWR _17196_/A sky130_fd_sc_hd__dfrtp_4
X_21549_ _17431_/Y _21549_/B VGND VGND VPWR VPWR _21549_/Y sky130_fd_sc_hd__nor2_4
X_15070_ _15193_/A _15070_/B _15070_/C _15069_/X VGND VGND VPWR VPWR _15070_/X sky130_fd_sc_hd__or4_4
X_12282_ _12220_/A _12282_/B _12282_/C _12281_/X VGND VGND VPWR VPWR _12283_/D sky130_fd_sc_hd__or4_4
XFILLER_126_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24268_ _24691_/CLK _17803_/X HRESETn VGND VGND VPWR VPWR _24268_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23234__A2 _22467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23069__C _23005_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14021_ _14003_/B _14016_/Y _14017_/Y _13995_/A _14020_/Y VGND VGND VPWR VPWR _14021_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_88_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23219_ _23219_/A _23310_/B VGND VGND VPWR VPWR _23219_/X sky130_fd_sc_hd__or2_4
X_24199_ _24305_/CLK _24199_/D HRESETn VGND VGND VPWR VPWR _24199_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22993__A1 _16485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16121__B1 _15962_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24339__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18760_ _18757_/B VGND VGND VPWR VPWR _18760_/Y sky130_fd_sc_hd__inv_2
X_15972_ _15966_/X _15969_/X _11809_/A _24748_/Q _15967_/X VGND VGND VPWR VPWR _15972_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_23_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17711_ _17708_/Y _17709_/Y _17710_/X VGND VGND VPWR VPWR _17711_/X sky130_fd_sc_hd__a21o_4
X_14923_ _25002_/Q _14922_/A _15064_/A _14922_/Y VGND VGND VPWR VPWR _14923_/X sky130_fd_sc_hd__o22a_4
X_18691_ _18758_/A _18757_/A _18626_/Y _18753_/C VGND VGND VPWR VPWR _18691_/X sky130_fd_sc_hd__or4_4
XFILLER_114_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17642_ _17642_/A _17642_/B _17641_/Y VGND VGND VPWR VPWR _17642_/X sky130_fd_sc_hd__and3_4
XFILLER_36_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14854_ _14845_/X _14853_/Y _24945_/Q _14845_/X VGND VGND VPWR VPWR _14854_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13805_ _13802_/Y _13796_/X _13803_/X _13804_/X VGND VGND VPWR VPWR _25260_/D sky130_fd_sc_hd__a2bb2o_4
X_17573_ _17573_/A VGND VGND VPWR VPWR _17662_/A sky130_fd_sc_hd__inv_2
X_11997_ _11990_/Y _11997_/B VGND VGND VPWR VPWR _11997_/Y sky130_fd_sc_hd__nor2_4
X_14785_ _14785_/A VGND VGND VPWR VPWR _17980_/A sky130_fd_sc_hd__inv_2
XFILLER_17_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19312_ _19311_/Y VGND VGND VPWR VPWR _19312_/X sky130_fd_sc_hd__buf_2
X_16524_ _16504_/A VGND VGND VPWR VPWR _16524_/X sky130_fd_sc_hd__buf_2
XANTENNA__15612__A _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23974__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13736_ _13735_/X VGND VGND VPWR VPWR _13736_/X sky130_fd_sc_hd__buf_2
XANTENNA__16188__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25198__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19243_ _19242_/X VGND VGND VPWR VPWR _19256_/A sky130_fd_sc_hd__inv_2
X_16455_ _16725_/A _16725_/B _22736_/A _21314_/B VGND VGND VPWR VPWR _16455_/X sky130_fd_sc_hd__and4_4
X_13667_ _20943_/A _24057_/Q _13667_/C _13666_/X VGND VGND VPWR VPWR _13667_/X sky130_fd_sc_hd__or4_4
XANTENNA__14228__A _25186_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15406_ _15406_/A _15390_/X VGND VGND VPWR VPWR _15406_/Y sky130_fd_sc_hd__nand2_4
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12618_ _12570_/Y _12565_/Y _12693_/B VGND VGND VPWR VPWR _12618_/X sky130_fd_sc_hd__or3_4
X_19174_ _14663_/D _19038_/B _19013_/X VGND VGND VPWR VPWR _19175_/A sky130_fd_sc_hd__or3_4
X_13598_ _11710_/A _13593_/X _13598_/C _14675_/C VGND VGND VPWR VPWR _13598_/X sky130_fd_sc_hd__or4_4
X_16386_ HWDATA[27] VGND VGND VPWR VPWR _16386_/X sky130_fd_sc_hd__buf_2
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18125_ _18054_/X _23816_/Q VGND VGND VPWR VPWR _18127_/B sky130_fd_sc_hd__or2_4
X_12549_ _24851_/Q VGND VGND VPWR VPWR _12549_/Y sky130_fd_sc_hd__inv_2
X_15337_ _15135_/Y _15344_/A VGND VGND VPWR VPWR _15338_/B sky130_fd_sc_hd__or2_4
XANTENNA__22681__B1 _22680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18056_ _18056_/A _18056_/B VGND VGND VPWR VPWR _18056_/X sky130_fd_sc_hd__or2_4
XANTENNA__24082__D _20952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15268_ _15250_/A _15267_/X _15174_/X VGND VGND VPWR VPWR _15268_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16360__B1 _16359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17007_ _17007_/A VGND VGND VPWR VPWR _17007_/Y sky130_fd_sc_hd__inv_2
X_14219_ _14219_/A VGND VGND VPWR VPWR _14220_/A sky130_fd_sc_hd__buf_2
XANTENNA__15059__A _15246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15199_ _15199_/A VGND VGND VPWR VPWR _15199_/X sky130_fd_sc_hd__buf_2
XFILLER_67_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24762__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15209__D _15171_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17274__A _17261_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25124__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18958_ _18957_/Y _18952_/X _16787_/X _18952_/X VGND VGND VPWR VPWR _23896_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24009__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25187__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17909_ _17909_/A VGND VGND VPWR VPWR _17909_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11814__A1_N _11811_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18889_ _18869_/X _18883_/X _23948_/Q _20974_/B _18886_/X VGND VGND VPWR VPWR _24109_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_67_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20920_ _16662_/Y _20814_/X _20845_/X _20919_/X VGND VGND VPWR VPWR _20920_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_8_235_0_HCLK clkbuf_8_235_0_HCLK/A VGND VGND VPWR VPWR _25356_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15769__A3 _15768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20851_ _20851_/A VGND VGND VPWR VPWR _20851_/Y sky130_fd_sc_hd__inv_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19365__B1 _19364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23570_ _23545_/CLK _23570_/D VGND VGND VPWR VPWR _19894_/A sky130_fd_sc_hd__dfxtp_4
X_20782_ _20781_/X VGND VGND VPWR VPWR _20782_/Y sky130_fd_sc_hd__inv_2
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22521_ _23327_/B VGND VGND VPWR VPWR _22522_/B sky130_fd_sc_hd__buf_2
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15926__B1 _12983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25240_ _24148_/CLK _25240_/D HRESETn VGND VGND VPWR VPWR _13851_/A sky130_fd_sc_hd__dfrtp_4
X_22452_ _12104_/Y _12060_/B _12014_/Y _13533_/B VGND VGND VPWR VPWR _22452_/X sky130_fd_sc_hd__o22a_4
X_21403_ _21403_/A _21395_/X _21402_/X VGND VGND VPWR VPWR _21403_/X sky130_fd_sc_hd__or3_4
XANTENNA__17449__A _24310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25171_ _24070_/CLK _25171_/D HRESETn VGND VGND VPWR VPWR _25171_/Q sky130_fd_sc_hd__dfrtp_4
X_22383_ _22383_/A _22301_/X _22383_/C _22383_/D VGND VGND VPWR VPWR _22383_/X sky130_fd_sc_hd__or4_4
X_24122_ _24117_/CLK _24122_/D HRESETn VGND VGND VPWR VPWR _18630_/A sky130_fd_sc_hd__dfrtp_4
X_21334_ _21334_/A _22172_/B VGND VGND VPWR VPWR _21334_/X sky130_fd_sc_hd__and2_4
XFILLER_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16351__B1 _16061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24326__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24053_ _24487_/CLK _24053_/D HRESETn VGND VGND VPWR VPWR _24053_/Q sky130_fd_sc_hd__dfrtp_4
X_21265_ _21498_/A _21263_/X _25258_/Q _21264_/X VGND VGND VPWR VPWR _21265_/X sky130_fd_sc_hd__o22a_4
XFILLER_46_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23004_ _23004_/A _22722_/B VGND VGND VPWR VPWR _23007_/B sky130_fd_sc_hd__or2_4
X_20216_ _20216_/A VGND VGND VPWR VPWR _20216_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21196_ _21196_/A _21196_/B _21196_/C VGND VGND VPWR VPWR _21196_/X sky130_fd_sc_hd__or3_4
XANTENNA__22090__A _22923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24432__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20147_ _19844_/X _13762_/X _19822_/C VGND VGND VPWR VPWR _20148_/A sky130_fd_sc_hd__or3_4
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_45_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20078_ _20095_/A VGND VGND VPWR VPWR _20078_/X sky130_fd_sc_hd__buf_2
X_24955_ _24955_/CLK _15448_/X HRESETn VGND VGND VPWR VPWR _13889_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_58_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13217__A _13162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11920_ _11916_/X VGND VGND VPWR VPWR _11920_/Y sky130_fd_sc_hd__inv_2
X_23906_ _23905_/CLK _23906_/D VGND VGND VPWR VPWR _13272_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24886_ _24889_/CLK _24886_/D HRESETn VGND VGND VPWR VPWR _24886_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16957__A2 _16955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11851_ HWDATA[3] VGND VGND VPWR VPWR _18254_/A sky130_fd_sc_hd__buf_2
XANTENNA__21434__A _23097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23837_ _25488_/CLK _19125_/X VGND VGND VPWR VPWR _19124_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16528__A _16528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14570_ _14570_/A _14570_/B VGND VGND VPWR VPWR _14571_/A sky130_fd_sc_hd__and2_4
XFILLER_60_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11782_ _11780_/Y _11777_/X _11781_/X _11777_/X VGND VGND VPWR VPWR _11782_/X sky130_fd_sc_hd__a2bb2o_4
X_23768_ _25503_/CLK _19323_/X VGND VGND VPWR VPWR _23768_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16262__A1_N _16261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17350__C _17350_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25291__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_HCLK clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13521_ _12026_/X VGND VGND VPWR VPWR _20953_/B sky130_fd_sc_hd__inv_2
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25507_ _24248_/CLK _11868_/X HRESETn VGND VGND VPWR VPWR _11864_/A sky130_fd_sc_hd__dfrtp_4
X_22719_ _22719_/A _22693_/Y _22711_/X _22718_/Y VGND VGND VPWR VPWR HRDATA[14] sky130_fd_sc_hd__or4_4
XFILLER_41_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23699_ _23683_/CLK _19519_/X VGND VGND VPWR VPWR _23699_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19108__B1 _19018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13452_ _13452_/A _19657_/A VGND VGND VPWR VPWR _13453_/C sky130_fd_sc_hd__or2_4
X_16240_ _22583_/A VGND VGND VPWR VPWR _16240_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25438_ _25425_/CLK _12446_/X HRESETn VGND VGND VPWR VPWR _12199_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22265__A _21570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12403_ _12385_/B _12391_/X _12402_/X _12398_/Y VGND VGND VPWR VPWR _12404_/A sky130_fd_sc_hd__a211o_4
X_13383_ _13297_/X _13375_/X _13383_/C VGND VGND VPWR VPWR _13383_/X sky130_fd_sc_hd__and3_4
X_16171_ _16169_/A VGND VGND VPWR VPWR _16172_/B sky130_fd_sc_hd__buf_2
X_25369_ _25356_/CLK _12930_/Y HRESETn VGND VGND VPWR VPWR _22706_/A sky130_fd_sc_hd__dfrtp_4
X_12334_ _24809_/Q VGND VGND VPWR VPWR _12334_/Y sky130_fd_sc_hd__inv_2
X_15122_ _15122_/A VGND VGND VPWR VPWR _15122_/Y sky130_fd_sc_hd__inv_2
X_15053_ _25021_/Q _15051_/Y _25015_/Q _15052_/Y VGND VGND VPWR VPWR _15054_/D sky130_fd_sc_hd__a2bb2o_4
X_19930_ _19930_/A VGND VGND VPWR VPWR _19943_/A sky130_fd_sc_hd__inv_2
Xclkbuf_7_127_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_255_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12265_ _12264_/X _24738_/Q _12280_/A _12231_/Y VGND VGND VPWR VPWR _12271_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14004_ _13997_/X _13998_/X _14001_/X _14040_/D VGND VGND VPWR VPWR _14042_/D sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_3_6_0_HCLK_A clkbuf_3_6_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19861_ _23582_/Q VGND VGND VPWR VPWR _19861_/Y sky130_fd_sc_hd__inv_2
X_12196_ _21065_/A VGND VGND VPWR VPWR _12196_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22430__A3 _22266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18812_ _18812_/A VGND VGND VPWR VPWR _18812_/Y sky130_fd_sc_hd__inv_2
X_19792_ _19792_/A VGND VGND VPWR VPWR _19792_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24102__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18743_ _18692_/A _18692_/B _18743_/C _18693_/A VGND VGND VPWR VPWR _18765_/B sky130_fd_sc_hd__or4_4
X_15955_ HWDATA[21] VGND VGND VPWR VPWR _15955_/X sky130_fd_sc_hd__buf_2
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14906_ _14903_/X _14904_/Y _25022_/Q _14905_/Y VGND VGND VPWR VPWR _14910_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17822__A _17758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18674_ _18603_/A VGND VGND VPWR VPWR _18674_/Y sky130_fd_sc_hd__inv_2
X_15886_ _15713_/A VGND VGND VPWR VPWR _15886_/X sky130_fd_sc_hd__buf_2
XFILLER_91_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25379__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17625_ _17557_/Y _17611_/B VGND VGND VPWR VPWR _17626_/B sky130_fd_sc_hd__or2_4
XFILLER_97_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14837_ _14825_/X _14836_/Y _14817_/C _14825_/X VGND VGND VPWR VPWR _25040_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18856__A2_N _18675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19347__B1 _19212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25308__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17556_ _24308_/Q VGND VGND VPWR VPWR _17585_/A sky130_fd_sc_hd__inv_2
XFILLER_63_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_65_0_HCLK clkbuf_8_65_0_HCLK/A VGND VGND VPWR VPWR _24077_/CLK sky130_fd_sc_hd__clkbuf_1
X_14768_ _14767_/X VGND VGND VPWR VPWR _14772_/B sky130_fd_sc_hd__inv_2
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16507_ _16506_/Y _16504_/X _16235_/X _16504_/X VGND VGND VPWR VPWR _16507_/X sky130_fd_sc_hd__a2bb2o_4
X_13719_ _13688_/B _13707_/X _13718_/Y _13714_/X _11667_/A VGND VGND VPWR VPWR _25275_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15908__B1 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17487_ _17486_/X VGND VGND VPWR VPWR _17487_/Y sky130_fd_sc_hd__inv_2
X_14699_ _21403_/A VGND VGND VPWR VPWR _21388_/A sky130_fd_sc_hd__inv_2
X_19226_ _13265_/B VGND VGND VPWR VPWR _19226_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16438_ _16436_/Y _16433_/X _16355_/X _16437_/X VGND VGND VPWR VPWR _16438_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13797__A _16355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19157_ _19157_/A VGND VGND VPWR VPWR _19157_/Y sky130_fd_sc_hd__inv_2
X_16369_ _12050_/X _15991_/B _15991_/C _16369_/D VGND VGND VPWR VPWR _16722_/A sky130_fd_sc_hd__or4_4
XFILLER_30_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18108_ _18204_/A _18108_/B VGND VGND VPWR VPWR _18108_/X sky130_fd_sc_hd__or2_4
X_19088_ _23851_/Q VGND VGND VPWR VPWR _19088_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16333__B1 _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18039_ _18224_/A _18039_/B _18039_/C VGND VGND VPWR VPWR _18040_/C sky130_fd_sc_hd__or3_4
XANTENNA__12851__D _12851_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21050_ _21024_/A VGND VGND VPWR VPWR _21050_/X sky130_fd_sc_hd__buf_2
XFILLER_114_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21519__A _24774_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20001_ _20000_/X VGND VGND VPWR VPWR _20014_/A sky130_fd_sc_hd__inv_2
XFILLER_114_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15517__A _15535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22709__A1 _24856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22185__A2 _22407_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21952_ _21952_/A _13815_/X VGND VGND VPWR VPWR _21952_/X sky130_fd_sc_hd__or2_4
X_24740_ _24792_/CLK _24740_/D HRESETn VGND VGND VPWR VPWR _22141_/A sky130_fd_sc_hd__dfrtp_4
X_20903_ _16673_/Y _20814_/X _20845_/X _20902_/Y VGND VGND VPWR VPWR _20904_/A sky130_fd_sc_hd__o22a_4
X_24671_ _24700_/CLK _16160_/X HRESETn VGND VGND VPWR VPWR _21691_/A sky130_fd_sc_hd__dfrtp_4
X_21883_ _21601_/A _21881_/X _21883_/C VGND VGND VPWR VPWR _21883_/X sky130_fd_sc_hd__and3_4
XANTENNA__25049__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23622_ _23388_/CLK _19746_/X VGND VGND VPWR VPWR _23622_/Q sky130_fd_sc_hd__dfxtp_4
X_20834_ _16709_/Y _20815_/X _20824_/X _20833_/Y VGND VGND VPWR VPWR _20834_/X sky130_fd_sc_hd__o22a_4
XFILLER_70_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14695__A1_N _21612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23553_ _24930_/CLK _19939_/X VGND VGND VPWR VPWR _19938_/A sky130_fd_sc_hd__dfxtp_4
X_20765_ _20765_/A VGND VGND VPWR VPWR _20765_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22893__B1 _24826_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22504_ _22504_/A VGND VGND VPWR VPWR _22504_/Y sky130_fd_sc_hd__inv_2
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21701__B _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23484_ _23467_/CLK _20129_/X VGND VGND VPWR VPWR _20125_/A sky130_fd_sc_hd__dfxtp_4
X_20696_ _15629_/Y _20677_/X _20686_/X _20695_/Y VGND VGND VPWR VPWR _20697_/A sky130_fd_sc_hd__o22a_4
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12189__B2 _24751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25223_ _23967_/CLK _14079_/X HRESETn VGND VGND VPWR VPWR _13990_/B sky130_fd_sc_hd__dfrtp_4
X_22435_ _22764_/A VGND VGND VPWR VPWR _22435_/X sky130_fd_sc_hd__buf_2
XFILLER_52_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22645__B1 _16042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19510__B1 _11955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24684__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25154_ _24102_/CLK _25154_/D HRESETn VGND VGND VPWR VPWR _18370_/B sky130_fd_sc_hd__dfstp_4
X_22366_ _22362_/X _22365_/X _14677_/X VGND VGND VPWR VPWR _22366_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_108_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24613__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24105_ _24322_/CLK _24105_/D HRESETn VGND VGND VPWR VPWR _20982_/A sky130_fd_sc_hd__dfrtp_4
X_21317_ _21325_/A VGND VGND VPWR VPWR _22885_/A sky130_fd_sc_hd__buf_2
X_25085_ _24376_/CLK _25085_/D HRESETn VGND VGND VPWR VPWR _25085_/Q sky130_fd_sc_hd__dfrtp_4
X_22297_ _16451_/A _22297_/B _22297_/C VGND VGND VPWR VPWR _22383_/A sky130_fd_sc_hd__and3_4
XFILLER_117_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16811__A _16807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22532__B _22727_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12050_ _12050_/A VGND VGND VPWR VPWR _12050_/X sky130_fd_sc_hd__buf_2
X_24036_ _24581_/CLK _24036_/D HRESETn VGND VGND VPWR VPWR _13659_/A sky130_fd_sc_hd__dfrtp_4
X_21248_ _21252_/A _19863_/Y VGND VGND VPWR VPWR _21248_/X sky130_fd_sc_hd__or2_4
XFILLER_85_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12343__A2_N _12341_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20333__A _20333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21179_ _21175_/X _21178_/X _24201_/Q VGND VGND VPWR VPWR _21180_/C sky130_fd_sc_hd__o21a_4
XFILLER_132_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19577__B1 _11955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15740_ _15740_/A VGND VGND VPWR VPWR _15740_/X sky130_fd_sc_hd__buf_2
X_12952_ _12944_/B _12944_/D VGND VGND VPWR VPWR _12955_/B sky130_fd_sc_hd__or2_4
XFILLER_58_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24938_ _24148_/CLK _15481_/X HRESETn VGND VGND VPWR VPWR _14881_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__25472__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11903_ _11874_/Y _11899_/Y _11886_/Y _11902_/X VGND VGND VPWR VPWR _11904_/A sky130_fd_sc_hd__a211o_4
XFILLER_2_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15671_ _15671_/A VGND VGND VPWR VPWR _22520_/A sky130_fd_sc_hd__buf_2
X_12883_ _12854_/B _12862_/X _12854_/A VGND VGND VPWR VPWR _12883_/X sky130_fd_sc_hd__o21a_4
X_24869_ _24847_/CLK _15722_/X HRESETn VGND VGND VPWR VPWR _12527_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_45_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25401__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17410_ _17387_/A _17401_/A _23984_/Q _20990_/B _17404_/A VGND VGND VPWR VPWR _24322_/D
+ sky130_fd_sc_hd__a32o_4
X_14622_ _14622_/A VGND VGND VPWR VPWR _14622_/Y sky130_fd_sc_hd__inv_2
X_11834_ _11831_/Y _11826_/X _11833_/X _11826_/X VGND VGND VPWR VPWR _11834_/X sky130_fd_sc_hd__a2bb2o_4
X_18390_ _21091_/A _17271_/X _18389_/Y VGND VGND VPWR VPWR _24177_/D sky130_fd_sc_hd__o21a_4
XFILLER_96_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21136__B1 _12054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17306_/X _17339_/X _17341_/C VGND VGND VPWR VPWR _24341_/D sky130_fd_sc_hd__and3_4
XFILLER_18_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21687__A1 _18272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11765_ _11763_/Y _11760_/X _11764_/X _11760_/X VGND VGND VPWR VPWR _11765_/X sky130_fd_sc_hd__a2bb2o_4
X_14553_ HREADY HSEL VGND VGND VPWR VPWR _14553_/Y sky130_fd_sc_hd__nand2_4
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _13503_/Y _13501_/X _11838_/X _13501_/X VGND VGND VPWR VPWR _25300_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17272_ _17235_/Y _17269_/X _17263_/B _17271_/X VGND VGND VPWR VPWR _17273_/A sky130_fd_sc_hd__a211o_4
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _13693_/C VGND VGND VPWR VPWR _13702_/A sky130_fd_sc_hd__inv_2
X_14484_ _14483_/Y _14481_/X _14391_/X _14481_/X VGND VGND VPWR VPWR _14484_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19011_ _19009_/Y _19005_/X _19010_/X _18988_/Y VGND VGND VPWR VPWR _23877_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16223_ _16223_/A VGND VGND VPWR VPWR _16223_/Y sky130_fd_sc_hd__inv_2
X_13435_ _13233_/A _13433_/X _13434_/X VGND VGND VPWR VPWR _13435_/X sky130_fd_sc_hd__and3_4
XANTENNA__13410__A _13156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13366_ _13366_/A _13366_/B _13365_/X VGND VGND VPWR VPWR _13366_/X sky130_fd_sc_hd__and3_4
X_16154_ _22144_/A VGND VGND VPWR VPWR _16154_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24354__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15105_ _15105_/A VGND VGND VPWR VPWR _15105_/Y sky130_fd_sc_hd__inv_2
X_12317_ _25330_/Q VGND VGND VPWR VPWR _12991_/B sky130_fd_sc_hd__inv_2
XFILLER_138_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13297_ _13177_/A VGND VGND VPWR VPWR _13297_/X sky130_fd_sc_hd__buf_2
X_16085_ _11739_/A _22493_/B VGND VGND VPWR VPWR _16086_/A sky130_fd_sc_hd__and2_4
XFILLER_108_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21984__D _21983_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12248_ _12248_/A VGND VGND VPWR VPWR _12248_/Y sky130_fd_sc_hd__inv_2
X_15036_ _15064_/A VGND VGND VPWR VPWR _15250_/A sky130_fd_sc_hd__buf_2
X_19913_ _23563_/Q VGND VGND VPWR VPWR _19913_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22403__A3 _21290_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11865__A HWDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19844_ _25267_/Q VGND VGND VPWR VPWR _19844_/X sky130_fd_sc_hd__buf_2
X_12179_ _25451_/Q VGND VGND VPWR VPWR _12179_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19775_ _19774_/X VGND VGND VPWR VPWR _19793_/A sky130_fd_sc_hd__inv_2
XANTENNA__16784__A1_N _15027_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16987_ _16987_/A VGND VGND VPWR VPWR _17034_/A sky130_fd_sc_hd__inv_2
X_18726_ _18658_/Y _18693_/X _18743_/C VGND VGND VPWR VPWR _18736_/A sky130_fd_sc_hd__or3_4
XFILLER_7_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15938_ _15937_/Y VGND VGND VPWR VPWR _15938_/X sky130_fd_sc_hd__buf_2
XFILLER_110_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18240__B1 _15747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18657_ _16557_/Y _24139_/Q _24522_/Q _18656_/Y VGND VGND VPWR VPWR _18660_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11863__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15869_ _15868_/X VGND VGND VPWR VPWR _15869_/X sky130_fd_sc_hd__buf_2
XFILLER_37_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25142__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17608_ _17582_/X _17600_/D _17560_/Y VGND VGND VPWR VPWR _17608_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15072__A _15187_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18588_ _18472_/A _18588_/B VGND VGND VPWR VPWR _18589_/B sky130_fd_sc_hd__or2_4
XANTENNA__21127__B1 _14377_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17539_ _24306_/Q VGND VGND VPWR VPWR _17559_/A sky130_fd_sc_hd__inv_2
XFILLER_127_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20550_ _14441_/Y _20533_/X _20547_/X _20549_/X VGND VGND VPWR VPWR _20551_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16554__B1 _16384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_9_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19209_ _19208_/Y _19203_/X _19117_/X _19203_/X VGND VGND VPWR VPWR _23808_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22627__B1 _24819_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20481_ _20488_/A _24073_/Q _20481_/C VGND VGND VPWR VPWR _20481_/X sky130_fd_sc_hd__and3_4
X_22220_ _22220_/A _19585_/A VGND VGND VPWR VPWR _22220_/X sky130_fd_sc_hd__and2_4
XANTENNA__20102__B2 _20095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24095__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22151_ _24439_/Q _21293_/X _22885_/A VGND VGND VPWR VPWR _22151_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24024__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21102_ _21826_/A VGND VGND VPWR VPWR _21103_/A sky130_fd_sc_hd__buf_2
XFILLER_133_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22082_ _14714_/X _22058_/Y _22066_/Y _22074_/Y _22081_/Y VGND VGND VPWR VPWR _22082_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_7_110_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_221_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21033_ _12604_/A _15654_/A _21031_/X _21032_/X VGND VGND VPWR VPWR _21034_/A sky130_fd_sc_hd__a211o_4
XANTENNA__12343__B2 _12345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18558__A _16448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23183__B _23182_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22984_ _22984_/A _22914_/B VGND VGND VPWR VPWR _22984_/X sky130_fd_sc_hd__and2_4
XFILLER_41_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24723_ _24345_/CLK _16025_/X HRESETn VGND VGND VPWR VPWR _24723_/Q sky130_fd_sc_hd__dfrtp_4
X_21935_ _21458_/A _21935_/B VGND VGND VPWR VPWR _21935_/X sky130_fd_sc_hd__or2_4
XANTENNA__11854__B1 _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21866_ _11720_/B VGND VGND VPWR VPWR _22425_/A sky130_fd_sc_hd__buf_2
X_24654_ _24654_/CLK _16215_/X HRESETn VGND VGND VPWR VPWR _24654_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16793__B1 _16720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _20816_/X VGND VGND VPWR VPWR _20909_/A sky130_fd_sc_hd__buf_2
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23605_ _23453_/CLK _23605_/D VGND VGND VPWR VPWR _23605_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19389__A _16786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22866__B1 _25525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21797_ _21452_/A _21795_/X _21796_/X VGND VGND VPWR VPWR _21797_/X sky130_fd_sc_hd__and3_4
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24585_ _24980_/CLK _24585_/D HRESETn VGND VGND VPWR VPWR _24585_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24865__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15710__A _15740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20748_ _20743_/X _20746_/Y _15599_/A _20747_/X VGND VGND VPWR VPWR _24012_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23536_ _23714_/CLK _23536_/D VGND VGND VPWR VPWR _19987_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23467_ _23467_/CLK _20173_/X VGND VGND VPWR VPWR _23467_/Q sky130_fd_sc_hd__dfxtp_4
X_20679_ _20678_/X VGND VGND VPWR VPWR _20770_/A sky130_fd_sc_hd__buf_2
XANTENNA__21150__C _21314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ _13269_/A _23377_/Q VGND VGND VPWR VPWR _13223_/B sky130_fd_sc_hd__or2_4
X_22418_ _22962_/A VGND VGND VPWR VPWR _22778_/A sky130_fd_sc_hd__buf_2
X_25206_ _25205_/CLK _14149_/X HRESETn VGND VGND VPWR VPWR _14116_/A sky130_fd_sc_hd__dfrtp_4
X_23398_ _23398_/CLK _20353_/X VGND VGND VPWR VPWR _20351_/A sky130_fd_sc_hd__dfxtp_4
X_13151_ _13212_/A VGND VGND VPWR VPWR _13248_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22349_ _21929_/A _19887_/Y _21191_/A VGND VGND VPWR VPWR _22349_/X sky130_fd_sc_hd__o21a_4
XFILLER_128_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25137_ _25137_/CLK _14392_/X HRESETn VGND VGND VPWR VPWR _20420_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_136_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12102_ _12119_/A VGND VGND VPWR VPWR _12102_/X sky130_fd_sc_hd__buf_2
XFILLER_124_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13082_ _12995_/A _13081_/X VGND VGND VPWR VPWR _13082_/X sky130_fd_sc_hd__or2_4
X_25068_ _25054_/CLK _14631_/X HRESETn VGND VGND VPWR VPWR _14613_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_3_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12033_ _12033_/A VGND VGND VPWR VPWR _12033_/Y sky130_fd_sc_hd__inv_2
X_16910_ _16105_/A _24269_/Q _16105_/Y _16909_/Y VGND VGND VPWR VPWR _16913_/C sky130_fd_sc_hd__o22a_4
XFILLER_105_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22397__A2 _22393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19798__B1 _19797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13531__B1 SCLK_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24019_ _24865_/CLK _20778_/X HRESETn VGND VGND VPWR VPWR _24019_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17890_ _24243_/Q VGND VGND VPWR VPWR _17900_/A sky130_fd_sc_hd__inv_2
XFILLER_137_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16841_ _14934_/Y _16837_/X _16600_/X _16840_/X VGND VGND VPWR VPWR _16841_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_5_15_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19560_ _18275_/X _20338_/B _19492_/X VGND VGND VPWR VPWR _19561_/A sky130_fd_sc_hd__or3_4
X_16772_ _15023_/Y _16770_/X _11821_/X _16770_/X VGND VGND VPWR VPWR _16772_/X sky130_fd_sc_hd__a2bb2o_4
X_13984_ _13984_/A _13980_/Y _13984_/C _13983_/X VGND VGND VPWR VPWR _13984_/X sky130_fd_sc_hd__and4_4
XFILLER_98_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18511_ _18460_/A _18514_/B _18487_/X VGND VGND VPWR VPWR _18511_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_46_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15723_ HWDATA[26] VGND VGND VPWR VPWR _15723_/X sky130_fd_sc_hd__buf_2
X_12935_ _22660_/A _12933_/A VGND VGND VPWR VPWR _12935_/X sky130_fd_sc_hd__or2_4
X_19491_ _17730_/X VGND VGND VPWR VPWR _20338_/A sky130_fd_sc_hd__buf_2
XFILLER_34_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18442_ _24167_/Q VGND VGND VPWR VPWR _18442_/Y sky130_fd_sc_hd__inv_2
X_15654_ _15654_/A VGND VGND VPWR VPWR _15655_/A sky130_fd_sc_hd__buf_2
X_12866_ _12882_/A VGND VGND VPWR VPWR _12866_/X sky130_fd_sc_hd__buf_2
XFILLER_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16784__B1 _16782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14605_ _14601_/B _14604_/Y _14599_/X _14602_/X _13582_/A VGND VGND VPWR VPWR _25074_/D
+ sky130_fd_sc_hd__a32o_4
X_11817_ HWDATA[11] VGND VGND VPWR VPWR _11818_/A sky130_fd_sc_hd__buf_2
X_18373_ _18369_/Y _18372_/X _24184_/Q _18372_/X VGND VGND VPWR VPWR _24185_/D sky130_fd_sc_hd__a2bb2o_4
X_15585_ _24901_/Q VGND VGND VPWR VPWR _22985_/A sky130_fd_sc_hd__inv_2
X_12797_ _25356_/Q _12795_/Y _25360_/Q _12796_/Y VGND VGND VPWR VPWR _12804_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19722__B1 _19721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17321_/B VGND VGND VPWR VPWR _17324_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15620__A _16057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14536_ _14018_/X VGND VGND VPWR VPWR _14536_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12270__B1 _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _25536_/Q VGND VGND VPWR VPWR _11748_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16536__B1 _16442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20238__A _20232_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24535__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_139_0_HCLK clkbuf_7_69_0_HCLK/X VGND VGND VPWR VPWR _23618_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17255_ _22659_/A _17249_/Y _17252_/X _17254_/X VGND VGND VPWR VPWR _17255_/X sky130_fd_sc_hd__or4_4
X_14467_ _14465_/Y _14466_/X _14395_/X _14466_/X VGND VGND VPWR VPWR _14467_/X sky130_fd_sc_hd__a2bb2o_4
X_11679_ _25278_/Q VGND VGND VPWR VPWR _13690_/A sky130_fd_sc_hd__inv_2
XFILLER_35_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16206_ _16204_/Y _16200_/X _15949_/X _16205_/X VGND VGND VPWR VPWR _24658_/D sky130_fd_sc_hd__a2bb2o_4
X_13418_ _13450_/A _13416_/X _13418_/C VGND VGND VPWR VPWR _13422_/B sky130_fd_sc_hd__and3_4
X_17186_ _23072_/A VGND VGND VPWR VPWR _17293_/A sky130_fd_sc_hd__inv_2
X_14398_ _14397_/Y _14394_/X _14239_/X _14384_/A VGND VGND VPWR VPWR _25135_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22624__A3 _22396_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16137_ _22595_/A VGND VGND VPWR VPWR _16137_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21832__A1 _14207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12573__B2 _24865_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13349_ _13413_/A _13349_/B _13349_/C VGND VGND VPWR VPWR _13350_/C sky130_fd_sc_hd__and3_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23268__B _23249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21069__A _21069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16068_ _16066_/Y _16060_/X _15471_/X _16067_/X VGND VGND VPWR VPWR _16068_/X sky130_fd_sc_hd__a2bb2o_4
X_15019_ _24446_/Q VGND VGND VPWR VPWR _15019_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23282__A1_N _12266_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25394__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22793__C1 _22510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21060__A2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19827_ _22212_/B _19824_/X _19780_/X _19824_/X VGND VGND VPWR VPWR _23595_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12803__A2_N _22708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15275__B1 _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25323__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17282__A _17260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12089__B1 _11862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19758_ HWDATA[5] VGND VGND VPWR VPWR _19758_/X sky130_fd_sc_hd__buf_2
XFILLER_37_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18709_ _18709_/A VGND VGND VPWR VPWR _18709_/Y sky130_fd_sc_hd__inv_2
X_19689_ _19689_/A VGND VGND VPWR VPWR _19689_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21720_ _21720_/A VGND VGND VPWR VPWR _21720_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16775__B1 _16604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21651_ _21459_/A _20035_/Y VGND VGND VPWR VPWR _21652_/C sky130_fd_sc_hd__or2_4
Xclkbuf_7_35_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_71_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22312__A2 _12096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20602_ _20602_/A VGND VGND VPWR VPWR _20602_/X sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_9_0_HCLK_A clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24370_ _24364_/CLK _24370_/D HRESETn VGND VGND VPWR VPWR _24370_/Q sky130_fd_sc_hd__dfrtp_4
X_21582_ _21582_/A _21582_/B VGND VGND VPWR VPWR _21582_/X sky130_fd_sc_hd__and2_4
XFILLER_127_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12261__B1 _12433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_98_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_98_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24276__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23321_ _24028_/Q _21278_/X _24060_/Q _21302_/X VGND VGND VPWR VPWR _23321_/Y sky130_fd_sc_hd__a22oi_4
X_20533_ _20556_/A VGND VGND VPWR VPWR _20533_/X sky130_fd_sc_hd__buf_2
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24205__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23252_ _20942_/Y _21581_/X _20803_/Y _22280_/A VGND VGND VPWR VPWR _23252_/X sky130_fd_sc_hd__o22a_4
X_20464_ _20488_/A VGND VGND VPWR VPWR _20485_/B sky130_fd_sc_hd__inv_2
XANTENNA__22319__A2_N _21549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23273__B1 _24872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22203_ _14749_/A _22199_/X _22202_/X VGND VGND VPWR VPWR _22203_/X sky130_fd_sc_hd__or3_4
XFILLER_106_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20087__B1 _20085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23183_ _23274_/A _23182_/X VGND VGND VPWR VPWR _23183_/X sky130_fd_sc_hd__and2_4
X_20395_ _20394_/X VGND VGND VPWR VPWR _20395_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_4_0_HCLK clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22134_ _24333_/Q _22646_/A _22792_/A VGND VGND VPWR VPWR _22134_/X sky130_fd_sc_hd__a21o_4
XFILLER_106_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22491__A1_N _17350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23025__B1 _12586_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13513__B1 _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22065_ _21763_/A _22062_/X _22064_/X VGND VGND VPWR VPWR _22065_/X sky130_fd_sc_hd__and3_4
XFILLER_0_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21016_ _21408_/A VGND VGND VPWR VPWR _21017_/B sky130_fd_sc_hd__buf_2
XFILLER_43_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25064__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15705__A _15713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21426__B _22998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11827__B1 _11825_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22967_ _22967_/A _22472_/B VGND VGND VPWR VPWR _22967_/X sky130_fd_sc_hd__or2_4
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12720_ _12595_/Y _12704_/X VGND VGND VPWR VPWR _12720_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__13225__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24706_ _24356_/CLK _16070_/X HRESETn VGND VGND VPWR VPWR _24706_/Q sky130_fd_sc_hd__dfrtp_4
X_21918_ _21663_/A VGND VGND VPWR VPWR _21944_/A sky130_fd_sc_hd__buf_2
XANTENNA__16766__B1 _15747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22898_ _21525_/A VGND VGND VPWR VPWR _22898_/X sky130_fd_sc_hd__buf_2
X_12651_ _12651_/A _12651_/B VGND VGND VPWR VPWR _12656_/B sky130_fd_sc_hd__or2_4
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24637_ _24643_/CLK _16262_/X HRESETn VGND VGND VPWR VPWR _24637_/Q sky130_fd_sc_hd__dfrtp_4
X_21849_ _21331_/X _21845_/X _21848_/X VGND VGND VPWR VPWR _21862_/B sky130_fd_sc_hd__o21ai_4
XFILLER_54_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ _24870_/Q VGND VGND VPWR VPWR _12582_/Y sky130_fd_sc_hd__inv_2
X_15370_ _15372_/A _15370_/B _15370_/C VGND VGND VPWR VPWR _24980_/D sky130_fd_sc_hd__and3_4
XFILLER_24_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24568_ _24435_/CLK _16444_/X HRESETn VGND VGND VPWR VPWR _15125_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_19_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14321_ _25159_/Q _14299_/Y _25158_/Q _14296_/B VGND VGND VPWR VPWR _14321_/X sky130_fd_sc_hd__o22a_4
XFILLER_129_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23519_ _23550_/CLK _20037_/X VGND VGND VPWR VPWR _20035_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__13598__C _13598_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24499_ _23434_/CLK _24499_/D HRESETn VGND VGND VPWR VPWR _13741_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ _24371_/Q VGND VGND VPWR VPWR _17041_/C sky130_fd_sc_hd__inv_2
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14252_ _23991_/Q _14248_/X _14251_/X VGND VGND VPWR VPWR _14252_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_7_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22273__A _22273_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13203_ _24190_/Q VGND VGND VPWR VPWR _13440_/A sky130_fd_sc_hd__buf_2
XFILLER_136_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14183_ _14173_/B _14181_/Y _14129_/X _14182_/Y _14132_/A VGND VGND VPWR VPWR _14184_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23999__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24647__CLK _24581_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13134_ _20779_/A _13120_/X _20761_/A VGND VGND VPWR VPWR _13135_/A sky130_fd_sc_hd__or3_4
X_18991_ _18991_/A VGND VGND VPWR VPWR _18991_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13504__B1 _11838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12307__B2 _24833_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13065_ _13052_/X VGND VGND VPWR VPWR _13065_/Y sky130_fd_sc_hd__inv_2
X_17942_ _17957_/A _17940_/X _17941_/X VGND VGND VPWR VPWR _17942_/X sky130_fd_sc_hd__and3_4
XFILLER_65_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12016_ _12019_/B VGND VGND VPWR VPWR _12016_/Y sky130_fd_sc_hd__inv_2
X_17873_ _24250_/Q _17872_/Y VGND VGND VPWR VPWR _17873_/X sky130_fd_sc_hd__or2_4
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15257__B1 _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18198__A _17995_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23319__A1 _22783_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20250__B1 _19771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16824_ _16801_/A VGND VGND VPWR VPWR _16840_/A sky130_fd_sc_hd__buf_2
X_19612_ _19612_/A VGND VGND VPWR VPWR _19612_/X sky130_fd_sc_hd__buf_2
XFILLER_78_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19543_ _23690_/Q VGND VGND VPWR VPWR _19543_/Y sky130_fd_sc_hd__inv_2
X_16755_ _24451_/Q VGND VGND VPWR VPWR _16755_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13967_ _13886_/X VGND VGND VPWR VPWR _13967_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22542__A2 _23226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15706_ _21154_/B VGND VGND VPWR VPWR _22123_/A sky130_fd_sc_hd__buf_2
XANTENNA__17830__A _17755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24787__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12918_ _12936_/A _12912_/X _12918_/C VGND VGND VPWR VPWR _12918_/X sky130_fd_sc_hd__and3_4
X_19474_ _22226_/B _19471_/X _11934_/X _19471_/X VGND VGND VPWR VPWR _19474_/X sky130_fd_sc_hd__a2bb2o_4
X_16686_ _16685_/Y _16683_/X _15745_/X _16683_/X VGND VGND VPWR VPWR _24480_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16757__B1 _16410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13898_ _13897_/X VGND VGND VPWR VPWR _13898_/Y sky130_fd_sc_hd__inv_2
X_18425_ _22809_/A _18540_/A _16256_/Y _18581_/A VGND VGND VPWR VPWR _18431_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21352__A _21352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24716__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15637_ _15636_/Y _15632_/X _14470_/X _15632_/X VGND VGND VPWR VPWR _24881_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12849_ _12849_/A _12849_/B _12849_/C _12849_/D VGND VGND VPWR VPWR _12849_/X sky130_fd_sc_hd__or4_4
XFILLER_76_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_2_0_HCLK_A clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18356_ _18363_/A _18353_/Y _18355_/Y VGND VGND VPWR VPWR _18356_/X sky130_fd_sc_hd__a21o_4
XANTENNA__12243__B1 _12430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15568_ _15563_/A VGND VGND VPWR VPWR _15568_/X sky130_fd_sc_hd__buf_2
XANTENNA__16509__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17307_ _22659_/A _17249_/Y _17346_/B _17247_/X VGND VGND VPWR VPWR _17307_/X sky130_fd_sc_hd__or4_4
X_14519_ _25095_/Q _14511_/X _25094_/Q _14513_/X VGND VGND VPWR VPWR _14519_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12794__B2 _24777_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18287_ _18287_/A VGND VGND VPWR VPWR _18287_/X sky130_fd_sc_hd__buf_2
X_15499_ _15490_/X VGND VGND VPWR VPWR _15499_/X sky130_fd_sc_hd__buf_2
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17238_ _17295_/A VGND VGND VPWR VPWR _17239_/A sky130_fd_sc_hd__inv_2
XANTENNA__12189__A2_N _24751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22183__A _22183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17169_ _17169_/A VGND VGND VPWR VPWR _17369_/A sky130_fd_sc_hd__buf_2
XANTENNA__16181__A _16180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20180_ _21765_/B _20175_/X _20092_/X _20175_/X VGND VGND VPWR VPWR _23464_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22911__A _21306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25504__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15496__B1 HADDR[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12214__A _22892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21569__B1 _21558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20241__B1 _15766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23870_ _23869_/CLK _23870_/D VGND VGND VPWR VPWR _19032_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16996__B1 _16044_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22821_ _22821_/A VGND VGND VPWR VPWR _22821_/X sky130_fd_sc_hd__buf_2
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25540_ _23384_/CLK _25540_/D HRESETn VGND VGND VPWR VPWR _11650_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16748__B1 _16398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22752_ _22751_/X VGND VGND VPWR VPWR _22752_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24457__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21703_ _21524_/X _21699_/Y _22705_/A _21702_/X VGND VGND VPWR VPWR _21703_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25471_ _25305_/CLK _12080_/X HRESETn VGND VGND VPWR VPWR _25471_/Q sky130_fd_sc_hd__dfrtp_4
X_22683_ _23126_/A VGND VGND VPWR VPWR _23056_/A sky130_fd_sc_hd__buf_2
XANTENNA__23089__A3 _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21634_ _21614_/X _21633_/X _21493_/X VGND VGND VPWR VPWR _21634_/Y sky130_fd_sc_hd__a21oi_4
X_24422_ _24427_/CLK _16817_/X HRESETn VGND VGND VPWR VPWR _24422_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21565_ _21559_/A _12054_/A VGND VGND VPWR VPWR _21565_/X sky130_fd_sc_hd__or2_4
XFILLER_21_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24353_ _24356_/CLK _24353_/D HRESETn VGND VGND VPWR VPWR _17295_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20516_ _20515_/X VGND VGND VPWR VPWR _20516_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_122_0_HCLK clkbuf_7_61_0_HCLK/X VGND VGND VPWR VPWR _24649_/CLK sky130_fd_sc_hd__clkbuf_1
X_23304_ _24803_/Q _23304_/B VGND VGND VPWR VPWR _23304_/X sky130_fd_sc_hd__or2_4
X_24284_ _24285_/CLK _17682_/X HRESETn VGND VGND VPWR VPWR _17494_/A sky130_fd_sc_hd__dfrtp_4
X_21496_ _24209_/Q _21264_/X VGND VGND VPWR VPWR _21496_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_185_0_HCLK clkbuf_7_92_0_HCLK/X VGND VGND VPWR VPWR _24309_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12537__B2 _12536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23235_ _22701_/A _23235_/B _23235_/C VGND VGND VPWR VPWR _23235_/X sky130_fd_sc_hd__and3_4
X_20447_ _20447_/A _20439_/X VGND VGND VPWR VPWR _20447_/X sky130_fd_sc_hd__and2_4
XANTENNA__18268__A3 _18267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20075__A3 _11867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23166_ _22879_/A VGND VGND VPWR VPWR _23166_/X sky130_fd_sc_hd__buf_2
X_20378_ _21163_/B _20373_/X _19885_/A _20360_/Y VGND VGND VPWR VPWR _23388_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22821__A _22821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25245__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22117_ _22111_/X _22113_/Y _22115_/Y _22116_/X _21547_/Y VGND VGND VPWR VPWR _22117_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_122_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23097_ _23097_/A VGND VGND VPWR VPWR _23097_/X sky130_fd_sc_hd__buf_2
XFILLER_0_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22048_ _22048_/A VGND VGND VPWR VPWR _22048_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21437__A _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14870_ _14870_/A _14870_/B VGND VGND VPWR VPWR _14871_/A sky130_fd_sc_hd__or2_4
XFILLER_85_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21980__B1 _21504_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13821_ _13821_/A VGND VGND VPWR VPWR _13822_/A sky130_fd_sc_hd__buf_2
XFILLER_112_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23999_ _24033_/CLK _20689_/Y HRESETn VGND VGND VPWR VPWR _23999_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12267__A1_N _12266_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16540_ _16539_/Y _16461_/A _16366_/X _16461_/A VGND VGND VPWR VPWR _24534_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24880__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13752_ _13752_/A VGND VGND VPWR VPWR _13752_/X sky130_fd_sc_hd__buf_2
XANTENNA__20535__A1 _14169_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22268__A _22407_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12703_ _12616_/B _12702_/X VGND VGND VPWR VPWR _12704_/B sky130_fd_sc_hd__or2_4
X_16471_ _24561_/Q VGND VGND VPWR VPWR _16471_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13683_ _11669_/Y _13683_/B VGND VGND VPWR VPWR _13684_/B sky130_fd_sc_hd__or2_4
XANTENNA__16266__A _14470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18210_ _17928_/A _18210_/B _18209_/X VGND VGND VPWR VPWR _18210_/X sky130_fd_sc_hd__and3_4
XANTENNA__24127__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15422_ _15422_/A _15421_/Y VGND VGND VPWR VPWR _15423_/B sky130_fd_sc_hd__or2_4
XFILLER_34_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12634_ _12636_/B VGND VGND VPWR VPWR _12635_/B sky130_fd_sc_hd__inv_2
X_19190_ _18189_/B VGND VGND VPWR VPWR _19190_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12225__B1 _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12776__A1 _25362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18141_ _14646_/X _18139_/X _18140_/X VGND VGND VPWR VPWR _18141_/X sky130_fd_sc_hd__and3_4
XFILLER_15_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15353_ _15298_/B _15352_/X VGND VGND VPWR VPWR _15354_/A sky130_fd_sc_hd__or2_4
XFILLER_12_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ _12565_/A VGND VGND VPWR VPWR _12565_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_81_0_HCLK clkbuf_7_81_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_81_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14304_ _14303_/X VGND VGND VPWR VPWR _14304_/Y sky130_fd_sc_hd__inv_2
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18072_ _18201_/A _18070_/X _18071_/X VGND VGND VPWR VPWR _18072_/X sky130_fd_sc_hd__and3_4
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23237__B1 _23172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15284_ _15246_/A _15278_/B _15283_/Y VGND VGND VPWR VPWR _24996_/D sky130_fd_sc_hd__and3_4
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12496_ _12278_/C _12469_/X _12412_/A _12494_/B VGND VGND VPWR VPWR _12496_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17809__B _17755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17023_ _24632_/Q VGND VGND VPWR VPWR _17023_/Y sky130_fd_sc_hd__inv_2
X_14235_ _25183_/Q VGND VGND VPWR VPWR _14235_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14166_ _14181_/B _14098_/X _14098_/D _14165_/X VGND VGND VPWR VPWR _14166_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18664__B1 _16613_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22460__B2 _22442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15478__B1 _15477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13117_ _13116_/X VGND VGND VPWR VPWR _25322_/D sky130_fd_sc_hd__inv_2
X_14097_ _14097_/A VGND VGND VPWR VPWR _14119_/C sky130_fd_sc_hd__inv_2
X_18974_ _23889_/Q VGND VGND VPWR VPWR _18974_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13048_ _13048_/A _13048_/B VGND VGND VPWR VPWR _13048_/X sky130_fd_sc_hd__or2_4
X_17925_ _17920_/A _17920_/B _15912_/X VGND VGND VPWR VPWR _17925_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24968__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17856_ _16918_/Y _17846_/X _17850_/X VGND VGND VPWR VPWR _17856_/X sky130_fd_sc_hd__or3_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16807_ _16807_/A VGND VGND VPWR VPWR _16807_/X sky130_fd_sc_hd__buf_2
XFILLER_94_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17787_ _17738_/X _17787_/B _17787_/C VGND VGND VPWR VPWR _24272_/D sky130_fd_sc_hd__and3_4
X_14999_ _14981_/X _16785_/A _14981_/X _16785_/A VGND VGND VPWR VPWR _14999_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16738_ _15015_/Y _16734_/X _16386_/X _16734_/X VGND VGND VPWR VPWR _16738_/X sky130_fd_sc_hd__a2bb2o_4
X_19526_ _21808_/B _19521_/X _11948_/X _19521_/X VGND VGND VPWR VPWR _19526_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24550__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19457_ _19456_/Y _19452_/X _19389_/X _19452_/X VGND VGND VPWR VPWR _19457_/X sky130_fd_sc_hd__a2bb2o_4
X_16669_ _22984_/A _16664_/X _16401_/X _16664_/X VGND VGND VPWR VPWR _24487_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18408_ _16249_/A _24153_/Q _16249_/Y _18469_/B VGND VGND VPWR VPWR _18408_/X sky130_fd_sc_hd__o22a_4
X_19388_ _18101_/B VGND VGND VPWR VPWR _19388_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22906__A _22186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18339_ _18338_/X VGND VGND VPWR VPWR _18340_/B sky130_fd_sc_hd__inv_2
XFILLER_37_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12209__A _25427_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21350_ _14190_/B _21350_/B VGND VGND VPWR VPWR _21547_/A sky130_fd_sc_hd__or2_4
X_20301_ _23418_/Q VGND VGND VPWR VPWR _22235_/B sky130_fd_sc_hd__inv_2
X_21281_ _15646_/A _15654_/A _21030_/A _21038_/B VGND VGND VPWR VPWR _21281_/X sky130_fd_sc_hd__or4_4
XANTENNA__18642__A1_N _16620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23020_ _14971_/A _22833_/X _22090_/X _23019_/X VGND VGND VPWR VPWR _23021_/C sky130_fd_sc_hd__a211o_4
X_20232_ _20232_/A VGND VGND VPWR VPWR _20232_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18655__B1 _24530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15469__B1 _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20163_ _23470_/Q VGND VGND VPWR VPWR _20163_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17735__A _17700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20094_ _20094_/A VGND VGND VPWR VPWR _20094_/Y sky130_fd_sc_hd__inv_2
X_24971_ _24980_/CLK _24971_/D HRESETn VGND VGND VPWR VPWR _24971_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23175__C _23174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12879__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22754__A2 _22821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11783__A _25526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19080__B1 _19056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23922_ _25219_/CLK _20531_/X HRESETn VGND VGND VPWR VPWR _23922_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16969__B1 _24730_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21407__D _21407_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24638__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23853_ _23854_/CLK _19082_/X VGND VGND VPWR VPWR _23853_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22804_ _24518_/Q _22523_/A _22524_/A _22803_/X VGND VGND VPWR VPWR _22805_/C sky130_fd_sc_hd__a211o_4
X_20996_ _20996_/A _20996_/B _23968_/Q VGND VGND VPWR VPWR _20996_/X sky130_fd_sc_hd__or3_4
X_23784_ _23847_/CLK _23784_/D VGND VGND VPWR VPWR _23784_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24291__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25523_ _24267_/CLK _25523_/D HRESETn VGND VGND VPWR VPWR _25523_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22735_ _16585_/A _21049_/X _21731_/X _22734_/X VGND VGND VPWR VPWR _22736_/C sky130_fd_sc_hd__a211o_4
XFILLER_53_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25454_ _24102_/CLK _12170_/X HRESETn VGND VGND VPWR VPWR SCLK_S3 sky130_fd_sc_hd__dfstp_4
XFILLER_55_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22666_ _16506_/Y _15854_/X VGND VGND VPWR VPWR _22666_/X sky130_fd_sc_hd__and2_4
X_24405_ _24407_/CLK _24405_/D HRESETn VGND VGND VPWR VPWR _24405_/Q sky130_fd_sc_hd__dfrtp_4
X_21617_ _21240_/X VGND VGND VPWR VPWR _21618_/A sky130_fd_sc_hd__buf_2
XFILLER_138_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25385_ _25385_/CLK _25385_/D HRESETn VGND VGND VPWR VPWR _12830_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12119__A _12119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22597_ _15609_/Y _22747_/B VGND VGND VPWR VPWR _22597_/X sky130_fd_sc_hd__and2_4
XANTENNA__25497__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12350_ _12349_/Y _24821_/Q _12349_/Y _24821_/Q VGND VGND VPWR VPWR _12350_/X sky130_fd_sc_hd__a2bb2o_4
X_24336_ _24334_/CLK _24336_/D HRESETn VGND VGND VPWR VPWR _17184_/A sky130_fd_sc_hd__dfrtp_4
X_21548_ _21548_/A _21548_/B VGND VGND VPWR VPWR _21548_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__25426__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12281_ _12263_/Y _12499_/A _12280_/Y VGND VGND VPWR VPWR _12281_/X sky130_fd_sc_hd__or3_4
X_21479_ _21484_/A _21479_/B VGND VGND VPWR VPWR _21480_/C sky130_fd_sc_hd__or2_4
X_24267_ _24267_/CLK _24267_/D HRESETn VGND VGND VPWR VPWR _24267_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14020_ _14018_/X _14020_/B VGND VGND VPWR VPWR _14020_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__18646__B1 _16590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23218_ _23217_/X VGND VGND VPWR VPWR _23218_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22551__A _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24198_ _24288_/CLK _24198_/D HRESETn VGND VGND VPWR VPWR _24198_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_134_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23149_ _23148_/X VGND VGND VPWR VPWR _23149_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15971_ _15966_/X _15969_/X _11803_/X _24749_/Q _15967_/X VGND VGND VPWR VPWR _24749_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_95_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17710_ _17707_/A _17713_/A VGND VGND VPWR VPWR _17710_/X sky130_fd_sc_hd__and2_4
XANTENNA__15880__B1 _11778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14922_ _14922_/A VGND VGND VPWR VPWR _14922_/Y sky130_fd_sc_hd__inv_2
X_18690_ _24129_/Q VGND VGND VPWR VPWR _18753_/C sky130_fd_sc_hd__inv_2
XANTENNA__20756__B2 _20747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20769__A1_N _20743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17641_ _17521_/Y _17641_/B VGND VGND VPWR VPWR _17641_/Y sky130_fd_sc_hd__nand2_4
XFILLER_64_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24379__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14853_ _14852_/X VGND VGND VPWR VPWR _14853_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24308__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13804_ _13795_/X VGND VGND VPWR VPWR _13804_/X sky130_fd_sc_hd__buf_2
XANTENNA__17380__A _17199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17572_ _17517_/Y _17676_/A _17512_/Y _17494_/Y VGND VGND VPWR VPWR _17572_/X sky130_fd_sc_hd__or4_4
XFILLER_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14784_ _25045_/Q _16880_/A _14783_/Y VGND VGND VPWR VPWR _25045_/D sky130_fd_sc_hd__o21a_4
XFILLER_63_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11996_ _11994_/A _11994_/B _11995_/Y VGND VGND VPWR VPWR _11997_/B sky130_fd_sc_hd__o21a_4
XANTENNA__21705__B1 _25358_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19311_ _19310_/X VGND VGND VPWR VPWR _19311_/Y sky130_fd_sc_hd__inv_2
X_16523_ _24540_/Q VGND VGND VPWR VPWR _16523_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13735_ _13735_/A VGND VGND VPWR VPWR _13735_/X sky130_fd_sc_hd__buf_2
X_19242_ _13755_/A _13752_/X _13735_/X _13762_/A VGND VGND VPWR VPWR _19242_/X sky130_fd_sc_hd__or4_4
XFILLER_32_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16454_ _16454_/A VGND VGND VPWR VPWR _21314_/B sky130_fd_sc_hd__inv_2
X_13666_ _24054_/Q _24053_/Q _13648_/X _20922_/B VGND VGND VPWR VPWR _13666_/X sky130_fd_sc_hd__or4_4
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15405_ _15384_/A _15392_/X _15404_/Y VGND VGND VPWR VPWR _24970_/D sky130_fd_sc_hd__and3_4
X_12617_ _12612_/X _12614_/X _12616_/X VGND VGND VPWR VPWR _12693_/B sky130_fd_sc_hd__or3_4
X_19173_ _19173_/A VGND VGND VPWR VPWR _19173_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13518__A1_N _13517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16385_ _15145_/Y _16382_/X _16384_/X _16382_/X VGND VGND VPWR VPWR _16385_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ _13815_/A _14433_/A VGND VGND VPWR VPWR _14675_/C sky130_fd_sc_hd__or2_4
XFILLER_34_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16724__A _23021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18124_ _18220_/A _18124_/B _18124_/C VGND VGND VPWR VPWR _18128_/B sky130_fd_sc_hd__and3_4
X_15336_ _15336_/A _15336_/B _15336_/C _15336_/D VGND VGND VPWR VPWR _15344_/A sky130_fd_sc_hd__or4_4
X_12548_ _25397_/Q VGND VGND VPWR VPWR _12708_/A sky130_fd_sc_hd__inv_2
XANTENNA__23943__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25167__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18055_ _18054_/X _19180_/A VGND VGND VPWR VPWR _18057_/B sky130_fd_sc_hd__or2_4
XFILLER_129_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15267_ _15267_/A _15267_/B VGND VGND VPWR VPWR _15267_/X sky130_fd_sc_hd__or2_4
XFILLER_32_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12479_ _12479_/A VGND VGND VPWR VPWR _25430_/D sky130_fd_sc_hd__inv_2
X_17006_ _16066_/Y _24364_/Q _24731_/Q _17005_/Y VGND VGND VPWR VPWR _17011_/B sky130_fd_sc_hd__a2bb2o_4
X_14218_ _25188_/Q VGND VGND VPWR VPWR _14218_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15198_ _15198_/A _15196_/X _15198_/C VGND VGND VPWR VPWR _15198_/X sky130_fd_sc_hd__and3_4
XANTENNA__22461__A _22786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_25_0_HCLK clkbuf_7_12_0_HCLK/X VGND VGND VPWR VPWR _25461_/CLK sky130_fd_sc_hd__clkbuf_1
X_14149_ _14146_/X _14148_/Y _25126_/Q _14146_/X VGND VGND VPWR VPWR _14149_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17555__A _17624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_88_0_HCLK clkbuf_8_89_0_HCLK/A VGND VGND VPWR VPWR _25029_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18957_ _18957_/A VGND VGND VPWR VPWR _18957_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15871__B1 _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17908_ _17895_/Y _17905_/A _17907_/X _17893_/A _17905_/Y VGND VGND VPWR VPWR _17908_/X
+ sky130_fd_sc_hd__a32o_4
X_18888_ _18869_/X _18883_/X _20974_/B _24110_/Q _18886_/X VGND VGND VPWR VPWR _18888_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24731__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17839_ _17841_/B VGND VGND VPWR VPWR _17840_/B sky130_fd_sc_hd__inv_2
XANTENNA__12849__D _12849_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24049__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20850_ _20850_/A VGND VGND VPWR VPWR _24036_/D sky130_fd_sc_hd__inv_2
XFILLER_130_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19509_ _23702_/Q VGND VGND VPWR VPWR _19509_/Y sky130_fd_sc_hd__inv_2
X_20781_ _15579_/Y _20676_/X _20706_/X _20780_/X VGND VGND VPWR VPWR _20781_/X sky130_fd_sc_hd__o22a_4
XFILLER_63_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14419__A _14408_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13323__A _13162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22520_ _22520_/A VGND VGND VPWR VPWR _23327_/B sky130_fd_sc_hd__buf_2
XANTENNA__15926__A1 _15655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22451_ _11686_/Y _21160_/X _13575_/Y _22505_/A VGND VGND VPWR VPWR _22451_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21402_ _21398_/X _21401_/X _14676_/X VGND VGND VPWR VPWR _21402_/X sky130_fd_sc_hd__o21a_4
X_22382_ _21821_/A _22381_/Y VGND VGND VPWR VPWR _22383_/D sky130_fd_sc_hd__nor2_4
X_25170_ _25461_/CLK _25170_/D HRESETn VGND VGND VPWR VPWR _25170_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22672__B2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21333_ _21333_/A VGND VGND VPWR VPWR _22172_/B sky130_fd_sc_hd__buf_2
XANTENNA__11778__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24121_ _24136_/CLK _18801_/Y HRESETn VGND VGND VPWR VPWR _24121_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21264_ _13791_/X VGND VGND VPWR VPWR _21264_/X sky130_fd_sc_hd__buf_2
XFILLER_135_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24052_ _24049_/CLK _24052_/D HRESETn VGND VGND VPWR VPWR _13664_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22371__A _21618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20215_ _20214_/Y _20212_/X _19755_/X _20212_/X VGND VGND VPWR VPWR _23451_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23003_ _22979_/X _22983_/X _22987_/Y _23002_/X VGND VGND VPWR VPWR HRDATA[21] sky130_fd_sc_hd__a211o_4
X_21195_ _21191_/X _21194_/X _24201_/Q VGND VGND VPWR VPWR _21196_/C sky130_fd_sc_hd__o21a_4
XFILLER_81_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20146_ _23476_/Q VGND VGND VPWR VPWR _20146_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24819__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19053__B1 _18961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20077_ _20077_/A VGND VGND VPWR VPWR _20095_/A sky130_fd_sc_hd__inv_2
XFILLER_58_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24954_ _24950_/CLK _24954_/D HRESETn VGND VGND VPWR VPWR _24954_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24472__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23905_ _23905_/CLK _23905_/D VGND VGND VPWR VPWR _13310_/B sky130_fd_sc_hd__dfxtp_4
X_24885_ _24885_/CLK _24885_/D HRESETn VGND VGND VPWR VPWR _15625_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24401__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15713__A _15713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11850_ _25510_/Q VGND VGND VPWR VPWR _11850_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23836_ _23884_/CLK _23836_/D VGND VGND VPWR VPWR _19126_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_45_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11781_ HWDATA[20] VGND VGND VPWR VPWR _11781_/X sky130_fd_sc_hd__buf_2
XANTENNA__17367__B1 _17271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23767_ _23660_/CLK _19326_/X VGND VGND VPWR VPWR _23767_/Q sky130_fd_sc_hd__dfxtp_4
X_20979_ _20979_/A VGND VGND VPWR VPWR _20979_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14329__A _14329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13520_ _20958_/B VGND VGND VPWR VPWR _20955_/B sky130_fd_sc_hd__buf_2
XANTENNA__13233__A _13233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21702__A3 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25506_ _25503_/CLK _25506_/D HRESETn VGND VGND VPWR VPWR _25506_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22718_ _22658_/A _22718_/B VGND VGND VPWR VPWR _22718_/Y sky130_fd_sc_hd__nor2_4
XFILLER_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22546__A _22546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12573__A2_N _24865_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23698_ _23682_/CLK _23698_/D VGND VGND VPWR VPWR _23698_/Q sky130_fd_sc_hd__dfxtp_4
X_13451_ _13246_/X _13451_/B VGND VGND VPWR VPWR _13451_/X sky130_fd_sc_hd__or2_4
XFILLER_9_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25437_ _25425_/CLK _12449_/X HRESETn VGND VGND VPWR VPWR _25437_/Q sky130_fd_sc_hd__dfrtp_4
X_22649_ _21064_/X _22649_/B VGND VGND VPWR VPWR _22649_/X sky130_fd_sc_hd__and2_4
X_12402_ _12410_/A VGND VGND VPWR VPWR _12402_/X sky130_fd_sc_hd__buf_2
X_16170_ RsRx_S0 _16169_/Y _14772_/B VGND VGND VPWR VPWR _16170_/X sky130_fd_sc_hd__a21o_4
X_13382_ _13314_/A _13378_/X _13382_/C VGND VGND VPWR VPWR _13383_/C sky130_fd_sc_hd__or3_4
X_25368_ _25368_/CLK _25368_/D HRESETn VGND VGND VPWR VPWR _25368_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25130__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25260__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15121_ _15121_/A _15121_/B _15121_/C _15120_/X VGND VGND VPWR VPWR _15121_/X sky130_fd_sc_hd__or4_4
X_12333_ _25324_/Q VGND VGND VPWR VPWR _13107_/A sky130_fd_sc_hd__inv_2
X_24319_ _24318_/CLK _24319_/D HRESETn VGND VGND VPWR VPWR _17420_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12588__A2_N _12586_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25299_ _25301_/CLK _25299_/D HRESETn VGND VGND VPWR VPWR _25299_/Q sky130_fd_sc_hd__dfrtp_4
X_15052_ _24453_/Q VGND VGND VPWR VPWR _15052_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22415__A1 _25362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12264_ _12263_/Y VGND VGND VPWR VPWR _12264_/X sky130_fd_sc_hd__buf_2
XFILLER_120_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_241_0_HCLK clkbuf_8_241_0_HCLK/A VGND VGND VPWR VPWR _24487_/CLK sky130_fd_sc_hd__clkbuf_1
X_14003_ _14003_/A _14003_/B _14003_/C _14002_/X VGND VGND VPWR VPWR _14040_/D sky130_fd_sc_hd__or4_4
X_12195_ _12284_/A _12193_/Y _25447_/Q _12194_/Y VGND VGND VPWR VPWR _12195_/X sky130_fd_sc_hd__a2bb2o_4
X_19860_ _19858_/Y _19859_/X _19794_/X _19859_/X VGND VGND VPWR VPWR _19860_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19292__B1 _19291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12511__A2_N _24853_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18811_ _18678_/Y _18784_/X _18724_/A _18809_/B VGND VGND VPWR VPWR _18812_/A sky130_fd_sc_hd__a211o_4
XFILLER_96_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19791_ _21748_/B _19784_/X _19790_/X _19784_/X VGND VGND VPWR VPWR _19791_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22179__B1 _22167_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15954_ _15938_/X VGND VGND VPWR VPWR _15954_/X sky130_fd_sc_hd__buf_2
X_18742_ _18742_/A VGND VGND VPWR VPWR _18759_/A sky130_fd_sc_hd__buf_2
X_14905_ _14905_/A VGND VGND VPWR VPWR _14905_/Y sky130_fd_sc_hd__inv_2
X_18673_ _18647_/X VGND VGND VPWR VPWR _18673_/Y sky130_fd_sc_hd__inv_2
X_15885_ _12792_/Y _15882_/X _11791_/X _15882_/X VGND VGND VPWR VPWR _24789_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24142__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15623__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14836_ _14810_/X _14834_/X _14231_/A _14835_/X VGND VGND VPWR VPWR _14836_/Y sky130_fd_sc_hd__a22oi_4
X_17624_ _17624_/A VGND VGND VPWR VPWR _17642_/A sky130_fd_sc_hd__buf_2
XFILLER_36_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17555_ _17624_/A VGND VGND VPWR VPWR _17617_/A sky130_fd_sc_hd__buf_2
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14767_ _16173_/A _14772_/A _14766_/X VGND VGND VPWR VPWR _14767_/X sky130_fd_sc_hd__or3_4
X_11979_ _11701_/B _11972_/X _11978_/Y VGND VGND VPWR VPWR _11979_/X sky130_fd_sc_hd__a21o_4
XANTENNA__14239__A _11862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16506_ _16506_/A VGND VGND VPWR VPWR _16506_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13718_ _13718_/A _13686_/X VGND VGND VPWR VPWR _13718_/Y sky130_fd_sc_hd__nand2_4
X_17486_ _24196_/Q _17468_/X _17484_/Y VGND VGND VPWR VPWR _17486_/X sky130_fd_sc_hd__o21a_4
X_14698_ _14686_/Y _14719_/A _14698_/C _14698_/D VGND VGND VPWR VPWR _14698_/X sky130_fd_sc_hd__or4_4
XFILLER_60_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16030__B1 _15962_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22456__A _21408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25348__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16437_ _16381_/A VGND VGND VPWR VPWR _16437_/X sky130_fd_sc_hd__buf_2
X_19225_ _19224_/Y _19222_/X _19133_/X _19222_/X VGND VGND VPWR VPWR _19225_/X sky130_fd_sc_hd__a2bb2o_4
X_13649_ _24046_/Q _24047_/Q _20889_/A _13649_/D VGND VGND VPWR VPWR _20900_/B sky130_fd_sc_hd__or4_4
XFILLER_38_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16454__A _16454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19156_ _19151_/Y _19154_/X _19155_/X _19154_/X VGND VGND VPWR VPWR _23828_/D sky130_fd_sc_hd__a2bb2o_4
X_16368_ _24598_/Q VGND VGND VPWR VPWR _16368_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18858__B1 _24561_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24093__D MSI_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17269__B _17261_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21510__D _21509_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18107_ _17982_/X _19412_/A VGND VGND VPWR VPWR _18109_/B sky130_fd_sc_hd__or2_4
Xclkbuf_6_51_0_HCLK clkbuf_6_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15319_ _15318_/X VGND VGND VPWR VPWR _24993_/D sky130_fd_sc_hd__inv_2
X_19087_ _22361_/B _19086_/X _16863_/X _19086_/X VGND VGND VPWR VPWR _19087_/X sky130_fd_sc_hd__a2bb2o_4
X_16299_ _24624_/Q VGND VGND VPWR VPWR _16299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17530__B1 _11811_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18038_ _18181_/A _18036_/X _18038_/C VGND VGND VPWR VPWR _18039_/C sky130_fd_sc_hd__and3_4
XFILLER_99_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20417__B1 _15647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22957__A2 _22513_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17285__A _17178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24983__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21519__B _21519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20000_ _17730_/X _18280_/X _20000_/C _18287_/X VGND VGND VPWR VPWR _20000_/X sky130_fd_sc_hd__or4_4
XANTENNA__16097__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24912__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19989_ _21804_/B _19982_/X _19988_/X _19982_/X VGND VGND VPWR VPWR _23536_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22709__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21951_ _21933_/X _21948_/X _21950_/X VGND VGND VPWR VPWR _21951_/X sky130_fd_sc_hd__a21o_4
XFILLER_95_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20902_ _13649_/D _20897_/X _20901_/Y VGND VGND VPWR VPWR _20902_/Y sky130_fd_sc_hd__a21oi_4
X_24670_ _24700_/CLK _24670_/D HRESETn VGND VGND VPWR VPWR _21513_/A sky130_fd_sc_hd__dfrtp_4
X_21882_ _21904_/A _21882_/B VGND VGND VPWR VPWR _21883_/C sky130_fd_sc_hd__or2_4
XFILLER_82_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _23388_/CLK _23621_/D VGND VGND VPWR VPWR _19747_/A sky130_fd_sc_hd__dfxtp_4
X_20833_ _13656_/A _13656_/B _20832_/Y VGND VGND VPWR VPWR _20833_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21145__A1 _14241_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21145__B2 _21355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23552_ _23711_/CLK _19941_/X VGND VGND VPWR VPWR _23552_/Q sky130_fd_sc_hd__dfxtp_4
X_20764_ _15590_/Y _20676_/X _20706_/X _20763_/Y VGND VGND VPWR VPWR _20765_/A sky130_fd_sc_hd__o22a_4
XFILLER_23_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25089__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22503_ _13813_/B _22501_/X _21587_/X _22502_/X VGND VGND VPWR VPWR _22504_/A sky130_fd_sc_hd__o22a_4
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20695_ _13126_/A _13126_/B _20694_/Y VGND VGND VPWR VPWR _20695_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23483_ _23467_/CLK _23483_/D VGND VGND VPWR VPWR _23483_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25018__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25222_ _25043_/CLK _14080_/X HRESETn VGND VGND VPWR VPWR _13990_/C sky130_fd_sc_hd__dfrtp_4
X_22434_ _22778_/A _22424_/Y _22428_/Y _22434_/D VGND VGND VPWR VPWR _22434_/X sky130_fd_sc_hd__or4_4
XANTENNA__22645__A1 _15709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22645__B2 _22915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25153_ _24109_/CLK _25153_/D HRESETn VGND VGND VPWR VPWR _25153_/Q sky130_fd_sc_hd__dfrtp_4
X_22365_ _21763_/A _22363_/X _22364_/X VGND VGND VPWR VPWR _22365_/X sky130_fd_sc_hd__and3_4
XFILLER_109_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24104_ _24612_/CLK _18896_/X HRESETn VGND VGND VPWR VPWR _20984_/A sky130_fd_sc_hd__dfrtp_4
X_21316_ _21316_/A VGND VGND VPWR VPWR _21325_/A sky130_fd_sc_hd__inv_2
X_22296_ _24509_/Q _21312_/X _22997_/A _22295_/X VGND VGND VPWR VPWR _22297_/C sky130_fd_sc_hd__a211o_4
X_25084_ _24376_/CLK _14578_/X HRESETn VGND VGND VPWR VPWR _25084_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20408__B1 _15766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21247_ _21247_/A _21245_/X _21247_/C VGND VGND VPWR VPWR _21247_/X sky130_fd_sc_hd__and3_4
XANTENNA__15708__A _15708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24035_ _24035_/CLK _24035_/D HRESETn VGND VGND VPWR VPWR _13658_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23070__A1 _24526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24653__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21178_ _24200_/Q _21176_/X _21178_/C VGND VGND VPWR VPWR _21178_/X sky130_fd_sc_hd__and3_4
XFILLER_77_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14638__A1 _14620_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_71_0_HCLK clkbuf_8_71_0_HCLK/A VGND VGND VPWR VPWR _25219_/CLK sky130_fd_sc_hd__clkbuf_1
X_20129_ _22370_/B _20128_/X _20079_/X _20128_/X VGND VGND VPWR VPWR _20129_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13228__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19026__B1 _18955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12951_ _12951_/A VGND VGND VPWR VPWR _25365_/D sky130_fd_sc_hd__inv_2
XFILLER_46_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24937_ _24957_/CLK _24937_/D HRESETn VGND VGND VPWR VPWR _24937_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11902_ RsRx_S1 _11902_/B VGND VGND VPWR VPWR _11902_/X sky130_fd_sc_hd__and2_4
X_15670_ _15670_/A VGND VGND VPWR VPWR _15671_/A sky130_fd_sc_hd__buf_2
X_12882_ _12882_/A VGND VGND VPWR VPWR _12884_/A sky130_fd_sc_hd__buf_2
X_24868_ _24868_/CLK _15724_/X HRESETn VGND VGND VPWR VPWR _24868_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16260__B1 _15471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14621_ _13638_/X _14620_/X VGND VGND VPWR VPWR _14622_/A sky130_fd_sc_hd__or2_4
X_11833_ _13835_/A VGND VGND VPWR VPWR _11833_/X sky130_fd_sc_hd__buf_2
X_23819_ _23818_/CLK _19179_/X VGND VGND VPWR VPWR _19178_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_33_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21136__A1 _12123_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _24780_/CLK _15873_/X HRESETn VGND VGND VPWR VPWR _23181_/A sky130_fd_sc_hd__dfrtp_4
X_17340_ _22659_/A _17337_/X VGND VGND VPWR VPWR _17341_/C sky130_fd_sc_hd__or2_4
XPHY_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14551_/X VGND VGND VPWR VPWR _23333_/A sky130_fd_sc_hd__buf_2
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ HWDATA[25] VGND VGND VPWR VPWR _11764_/X sky130_fd_sc_hd__buf_2
XANTENNA__12821__B1 _25383_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25441__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _25300_/Q VGND VGND VPWR VPWR _13503_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17279_/A VGND VGND VPWR VPWR _17271_/X sky130_fd_sc_hd__buf_2
X_14483_ _14483_/A VGND VGND VPWR VPWR _14483_/Y sky130_fd_sc_hd__inv_2
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _25270_/Q _24215_/Q _13729_/A _11694_/Y VGND VGND VPWR VPWR _11695_/X sky130_fd_sc_hd__o22a_4
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19010_ _17442_/X VGND VGND VPWR VPWR _19010_/X sky130_fd_sc_hd__buf_2
XFILLER_109_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16222_ _16221_/Y _16217_/X _15964_/X _16217_/X VGND VGND VPWR VPWR _24651_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13434_ _13248_/A _19124_/A VGND VGND VPWR VPWR _13434_/X sky130_fd_sc_hd__or2_4
X_16153_ _16151_/Y _16152_/X _16061_/X _16152_/X VGND VGND VPWR VPWR _16153_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19501__B2 _19500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13365_ _13461_/A _13365_/B _13364_/X VGND VGND VPWR VPWR _13365_/X sky130_fd_sc_hd__or3_4
XFILLER_6_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15104_ _24970_/Q VGND VGND VPWR VPWR _15392_/A sky130_fd_sc_hd__inv_2
X_12316_ _12314_/A _24826_/Q _12988_/A _12315_/Y VGND VGND VPWR VPWR _12326_/A sky130_fd_sc_hd__o22a_4
X_16084_ _15854_/X VGND VGND VPWR VPWR _22493_/B sky130_fd_sc_hd__buf_2
X_13296_ _13198_/X _13295_/X _25318_/Q _13258_/X VGND VGND VPWR VPWR _13296_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15035_ _14926_/X _24452_/Q _14926_/X _24452_/Q VGND VGND VPWR VPWR _15035_/X sky130_fd_sc_hd__a2bb2o_4
X_19912_ _19908_/Y _19911_/X _19777_/X _19911_/X VGND VGND VPWR VPWR _23564_/D sky130_fd_sc_hd__a2bb2o_4
X_12247_ _12286_/B _24752_/Q _12284_/A _12193_/Y VGND VGND VPWR VPWR _12251_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24394__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19843_ _23588_/Q VGND VGND VPWR VPWR _19843_/Y sky130_fd_sc_hd__inv_2
X_12178_ _12475_/A _24746_/Q _12475_/A _24746_/Q VGND VGND VPWR VPWR _12178_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19774_ _13736_/X _13762_/X _19845_/C VGND VGND VPWR VPWR _19774_/X sky130_fd_sc_hd__or3_4
X_16986_ _24705_/Q _16985_/A _16071_/Y _16985_/Y VGND VGND VPWR VPWR _16989_/C sky130_fd_sc_hd__o22a_4
X_18725_ _18725_/A VGND VGND VPWR VPWR _18725_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21355__A _21355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15937_ _15967_/A VGND VGND VPWR VPWR _15937_/Y sky130_fd_sc_hd__inv_2
X_15868_ _15900_/A VGND VGND VPWR VPWR _15868_/X sky130_fd_sc_hd__buf_2
X_18656_ _24133_/Q VGND VGND VPWR VPWR _18656_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25529__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14819_ _14819_/A _14819_/B _14819_/C VGND VGND VPWR VPWR _14819_/X sky130_fd_sc_hd__and3_4
X_17607_ _17617_/A _17607_/B _17606_/X VGND VGND VPWR VPWR _24305_/D sky130_fd_sc_hd__and3_4
X_15799_ _15809_/A VGND VGND VPWR VPWR _15799_/X sky130_fd_sc_hd__buf_2
X_18587_ _18472_/A _18588_/B VGND VGND VPWR VPWR _18589_/A sky130_fd_sc_hd__nand2_4
XFILLER_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22324__B1 _22311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17538_ _11773_/Y _17543_/A _25517_/Q _17499_/Y VGND VGND VPWR VPWR _17538_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22186__A _22186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17469_ _17466_/Y _17467_/Y _17468_/X VGND VGND VPWR VPWR _17469_/X sky130_fd_sc_hd__a21o_4
XANTENNA__25111__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19208_ _19208_/A VGND VGND VPWR VPWR _19208_/Y sky130_fd_sc_hd__inv_2
X_20480_ _20487_/A _20479_/X VGND VGND VPWR VPWR _20480_/X sky130_fd_sc_hd__or2_4
XANTENNA__22627__A1 _22476_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22627__B2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19139_ _19139_/A VGND VGND VPWR VPWR _19139_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17503__B1 _11756_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22150_ _15077_/A _22927_/A VGND VGND VPWR VPWR _22153_/B sky130_fd_sc_hd__or2_4
XFILLER_69_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21101_ _23997_/Q VGND VGND VPWR VPWR _21101_/Y sky130_fd_sc_hd__inv_2
X_22081_ _21767_/X _22080_/X _14714_/X VGND VGND VPWR VPWR _22081_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__15528__A _24919_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14432__A _25124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21032_ _21006_/B _21074_/B VGND VGND VPWR VPWR _21032_/X sky130_fd_sc_hd__and2_4
XANTENNA__15247__B _15171_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_58_0_HCLK clkbuf_7_58_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19008__B1 _18940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22983_ _22981_/X _22982_/X _23117_/C VGND VGND VPWR VPWR _22983_/X sky130_fd_sc_hd__or3_4
XFILLER_95_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16359__A _16359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22563__B1 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11791__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24722_ _24712_/CLK _16028_/X HRESETn VGND VGND VPWR VPWR _24722_/Q sky130_fd_sc_hd__dfrtp_4
X_21934_ _21455_/A _21934_/B VGND VGND VPWR VPWR _21934_/X sky130_fd_sc_hd__or2_4
XFILLER_41_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15045__B2 _24447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24653_ _24162_/CLK _16218_/X HRESETn VGND VGND VPWR VPWR _16216_/A sky130_fd_sc_hd__dfrtp_4
X_21865_ _24776_/Q _21863_/X _23005_/C _24846_/Q _21067_/A VGND VGND VPWR VPWR _21865_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _23660_/CLK _19804_/X VGND VGND VPWR VPWR _13171_/B sky130_fd_sc_hd__dfxtp_4
X_20816_ _20812_/Y _13669_/Y VGND VGND VPWR VPWR _20816_/X sky130_fd_sc_hd__or2_4
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24584_ _24980_/CLK _24584_/D HRESETn VGND VGND VPWR VPWR _15122_/A sky130_fd_sc_hd__dfrtp_4
X_21796_ _21658_/A _21796_/B VGND VGND VPWR VPWR _21796_/X sky130_fd_sc_hd__or2_4
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23535_ _23533_/CLK _23535_/D VGND VGND VPWR VPWR _23535_/Q sky130_fd_sc_hd__dfxtp_4
X_20747_ _20747_/A VGND VGND VPWR VPWR _20747_/X sky130_fd_sc_hd__buf_2
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16094__A _16094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23466_ _23562_/CLK _23466_/D VGND VGND VPWR VPWR _20174_/A sky130_fd_sc_hd__dfxtp_4
X_20678_ _20674_/Y _13139_/Y VGND VGND VPWR VPWR _20678_/X sky130_fd_sc_hd__or2_4
XFILLER_104_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25205_ _25205_/CLK _14152_/X HRESETn VGND VGND VPWR VPWR _25205_/Q sky130_fd_sc_hd__dfrtp_4
X_22417_ _22383_/X _22399_/X _22417_/C _22417_/D VGND VGND VPWR VPWR HRDATA[7] sky130_fd_sc_hd__or4_4
XFILLER_104_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23397_ _23398_/CLK _20355_/X VGND VGND VPWR VPWR _20354_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_100_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13150_ _24190_/Q VGND VGND VPWR VPWR _13212_/A sky130_fd_sc_hd__inv_2
XANTENNA__24834__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25136_ _25178_/CLK _14396_/X HRESETn VGND VGND VPWR VPWR _14393_/A sky130_fd_sc_hd__dfrtp_4
X_22348_ _21945_/A _22348_/B VGND VGND VPWR VPWR _22348_/X sky130_fd_sc_hd__or2_4
X_12101_ _12101_/A VGND VGND VPWR VPWR _12119_/A sky130_fd_sc_hd__inv_2
XFILLER_30_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13081_ _12363_/Y _13081_/B VGND VGND VPWR VPWR _13081_/X sky130_fd_sc_hd__or2_4
X_25067_ _25054_/CLK _25067_/D HRESETn VGND VGND VPWR VPWR _21958_/A sky130_fd_sc_hd__dfrtp_4
X_22279_ _16704_/Y _22406_/B VGND VGND VPWR VPWR _22279_/X sky130_fd_sc_hd__and2_4
XFILLER_78_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12032_ _12031_/Y _12029_/X _12033_/A _12029_/X VGND VGND VPWR VPWR _25481_/D sky130_fd_sc_hd__a2bb2o_4
X_24018_ _24018_/CLK _20775_/X HRESETn VGND VGND VPWR VPWR _13120_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15808__B1 _11774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16840_ _16840_/A VGND VGND VPWR VPWR _16840_/X sky130_fd_sc_hd__buf_2
X_16771_ _16769_/Y _16770_/X _15752_/X _16770_/X VGND VGND VPWR VPWR _16771_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15823__A3 _15750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13983_ _13983_/A VGND VGND VPWR VPWR _13983_/X sky130_fd_sc_hd__buf_2
XFILLER_24_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22554__B1 _24713_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15722_ _12527_/Y _15718_/X _11757_/X _15721_/X VGND VGND VPWR VPWR _15722_/X sky130_fd_sc_hd__a2bb2o_4
X_18510_ _18460_/B _18517_/B VGND VGND VPWR VPWR _18514_/B sky130_fd_sc_hd__or2_4
X_12934_ _25368_/Q _12933_/Y VGND VGND VPWR VPWR _12934_/X sky130_fd_sc_hd__or2_4
X_19490_ _23708_/Q VGND VGND VPWR VPWR _22325_/B sky130_fd_sc_hd__inv_2
XANTENNA__16233__B1 _16231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15653_ _15653_/A VGND VGND VPWR VPWR _15654_/A sky130_fd_sc_hd__inv_2
X_18441_ _16199_/Y _24171_/Q _24654_/Q _18524_/A VGND VGND VPWR VPWR _18444_/C sky130_fd_sc_hd__a2bb2o_4
X_12865_ _12838_/A VGND VGND VPWR VPWR _12882_/A sky130_fd_sc_hd__inv_2
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14604_ _13582_/Y _14563_/B VGND VGND VPWR VPWR _14604_/Y sky130_fd_sc_hd__nand2_4
X_11816_ _11794_/X VGND VGND VPWR VPWR _11816_/X sky130_fd_sc_hd__buf_2
X_18372_ _18377_/A VGND VGND VPWR VPWR _18372_/X sky130_fd_sc_hd__buf_2
X_15584_ _15583_/Y _15581_/X _11774_/X _15581_/X VGND VGND VPWR VPWR _24902_/D sky130_fd_sc_hd__a2bb2o_4
X_12796_ _24777_/Q VGND VGND VPWR VPWR _12796_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17306_/X _17323_/B _17322_/Y VGND VGND VPWR VPWR _24346_/D sky130_fd_sc_hd__and3_4
XPHY_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _20531_/A VGND VGND VPWR VPWR _14535_/Y sky130_fd_sc_hd__inv_2
XPHY_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11745_/Y _11742_/X _11746_/X _11742_/X VGND VGND VPWR VPWR _11747_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12270__B2 _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17254_ _17254_/A _17203_/Y _17254_/C _17253_/Y VGND VGND VPWR VPWR _17254_/X sky130_fd_sc_hd__or4_4
XANTENNA__22609__A1 _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ _14453_/Y VGND VGND VPWR VPWR _14466_/X sky130_fd_sc_hd__buf_2
XFILLER_30_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _25273_/Q _11677_/A _13685_/A _11677_/Y VGND VGND VPWR VPWR _11678_/X sky130_fd_sc_hd__o22a_4
X_16205_ _16217_/A VGND VGND VPWR VPWR _16205_/X sky130_fd_sc_hd__buf_2
X_13417_ _13417_/A _19699_/A VGND VGND VPWR VPWR _13418_/C sky130_fd_sc_hd__or2_4
X_17185_ _16345_/A _17184_/A _16345_/Y _17246_/B VGND VGND VPWR VPWR _17191_/B sky130_fd_sc_hd__o22a_4
XANTENNA__19486__B1 _11955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22085__A2 _21073_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14397_ _25135_/Q VGND VGND VPWR VPWR _14397_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16136_ _16135_/Y _16131_/X _11813_/X _16131_/X VGND VGND VPWR VPWR _16136_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24575__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13348_ _13312_/A _13348_/B VGND VGND VPWR VPWR _13349_/C sky130_fd_sc_hd__or2_4
XFILLER_6_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24504__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16067_ _15995_/X VGND VGND VPWR VPWR _16067_/X sky130_fd_sc_hd__buf_2
XANTENNA__19238__B1 _19191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13279_ _13317_/A _19689_/A VGND VGND VPWR VPWR _13280_/C sky130_fd_sc_hd__or2_4
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15018_ _25025_/Q _24463_/Q _15166_/C _15017_/Y VGND VGND VPWR VPWR _15021_/C sky130_fd_sc_hd__o22a_4
XANTENNA__12325__A2 _24814_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19826_ _23595_/Q VGND VGND VPWR VPWR _22212_/B sky130_fd_sc_hd__inv_2
XFILLER_96_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16472__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19757_ _19757_/A VGND VGND VPWR VPWR _19757_/Y sky130_fd_sc_hd__inv_2
X_16969_ _24724_/Q _17035_/A _24730_/Q _17025_/B VGND VGND VPWR VPWR _16971_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18708_ _18698_/C _18705_/X _18701_/B _18707_/X VGND VGND VPWR VPWR _18709_/A sky130_fd_sc_hd__a211o_4
X_19688_ _19687_/Y _19685_/X _19642_/X _19685_/X VGND VGND VPWR VPWR _19688_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25363__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20020__B2 _20014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18639_ _24114_/Q VGND VGND VPWR VPWR _18639_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22628__B _22592_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21650_ _21650_/A _21650_/B VGND VGND VPWR VPWR _21652_/B sky130_fd_sc_hd__or2_4
XFILLER_33_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20601_ _20601_/A _20495_/X VGND VGND VPWR VPWR _20601_/X sky130_fd_sc_hd__and2_4
X_21581_ _22824_/A VGND VGND VPWR VPWR _21581_/X sky130_fd_sc_hd__buf_2
XFILLER_123_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23320_ _22782_/A _23320_/B VGND VGND VPWR VPWR _23320_/Y sky130_fd_sc_hd__nor2_4
X_20532_ _20562_/A VGND VGND VPWR VPWR _20556_/A sky130_fd_sc_hd__inv_2
XFILLER_137_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22644__A _24612_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20463_ _20443_/B _20601_/A _14541_/A _20425_/X VGND VGND VPWR VPWR _24076_/D sky130_fd_sc_hd__a211o_4
XANTENNA__23273__A1 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23251_ _12385_/A _22489_/X _23250_/X VGND VGND VPWR VPWR _23251_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_118_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22202_ _22078_/X _22202_/B _22201_/X VGND VGND VPWR VPWR _22202_/X sky130_fd_sc_hd__and3_4
Xclkbuf_5_21_0_HCLK clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20394_ _20978_/B _14096_/C VGND VGND VPWR VPWR _20394_/X sky130_fd_sc_hd__or2_4
X_23182_ _23034_/X _23181_/X _22968_/X _12527_/A _23102_/X VGND VGND VPWR VPWR _23182_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__11772__B1 _11771_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24245__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22133_ _21098_/A VGND VGND VPWR VPWR _22646_/A sky130_fd_sc_hd__buf_2
XFILLER_121_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12316__A2 _24826_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22064_ _22068_/A _20110_/Y VGND VGND VPWR VPWR _22064_/X sky130_fd_sc_hd__or2_4
XFILLER_82_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21015_ _21015_/A VGND VGND VPWR VPWR _21408_/A sky130_fd_sc_hd__buf_2
XFILLER_134_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23194__B _23226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23328__A2 _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15805__A3 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22000__A2 _22727_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_145_0_HCLK clkbuf_7_72_0_HCLK/X VGND VGND VPWR VPWR _24214_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_56_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22966_ _23143_/A _22966_/B VGND VGND VPWR VPWR _22979_/B sky130_fd_sc_hd__and2_4
XANTENNA__16215__B1 _15957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22819__A _21275_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24705_ _24356_/CLK _16072_/X HRESETn VGND VGND VPWR VPWR _24705_/Q sky130_fd_sc_hd__dfrtp_4
X_21917_ _21191_/A VGND VGND VPWR VPWR _21917_/X sky130_fd_sc_hd__buf_2
XANTENNA__21723__A _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22897_ _22897_/A _22897_/B VGND VGND VPWR VPWR _22905_/C sky130_fd_sc_hd__and2_4
XFILLER_82_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25033__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12650_ _12665_/A _12618_/X _12620_/B _12611_/X VGND VGND VPWR VPWR _12651_/B sky130_fd_sc_hd__or4_4
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24636_ _24643_/CLK _24636_/D HRESETn VGND VGND VPWR VPWR _24636_/Q sky130_fd_sc_hd__dfrtp_4
X_21848_ _21566_/X _21846_/X _21560_/X _21847_/X VGND VGND VPWR VPWR _21848_/X sky130_fd_sc_hd__o22a_4
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ _25392_/Q VGND VGND VPWR VPWR _12616_/B sky130_fd_sc_hd__inv_2
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24567_ _24435_/CLK _24567_/D HRESETn VGND VGND VPWR VPWR _16445_/A sky130_fd_sc_hd__dfrtp_4
X_21779_ _21636_/X _21778_/X _13799_/A _18261_/A VGND VGND VPWR VPWR _21779_/X sky130_fd_sc_hd__o22a_4
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14320_ _14305_/Y _14319_/X _13488_/A _14311_/X VGND VGND VPWR VPWR _25160_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13241__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14529__B1 _25103_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23518_ _23550_/CLK _20039_/X VGND VGND VPWR VPWR _20038_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_12_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24498_ _23498_/CLK _24498_/D HRESETn VGND VGND VPWR VPWR _16630_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ _14251_/A _14244_/X _15428_/A _14251_/D VGND VGND VPWR VPWR _14251_/X sky130_fd_sc_hd__or4_4
XFILLER_8_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17648__A _17565_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23449_ _23660_/CLK _23449_/D VGND VGND VPWR VPWR _23449_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22273__B _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13202_ _24191_/Q VGND VGND VPWR VPWR _13413_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14182_ _14182_/A VGND VGND VPWR VPWR _14182_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13133_ _13133_/A _13133_/B _24012_/Q _20740_/A VGND VGND VPWR VPWR _20761_/A sky130_fd_sc_hd__or4_4
XANTENNA__23016__A1 _21409_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25119_ _25101_/CLK _25119_/D HRESETn VGND VGND VPWR VPWR _25119_/Q sky130_fd_sc_hd__dfstp_4
X_18990_ _18986_/Y _18989_/X _17418_/X _18989_/X VGND VGND VPWR VPWR _23884_/D sky130_fd_sc_hd__a2bb2o_4
X_13064_ _13049_/A _13064_/B _13063_/Y VGND VGND VPWR VPWR _25338_/D sky130_fd_sc_hd__and3_4
X_17941_ _17956_/A _19195_/A VGND VGND VPWR VPWR _17941_/X sky130_fd_sc_hd__or2_4
XANTENNA__19582__B _21143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12015_ _12015_/A _11994_/X VGND VGND VPWR VPWR _12019_/B sky130_fd_sc_hd__and2_4
X_17872_ _17850_/D VGND VGND VPWR VPWR _17872_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19640__B1 _19426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16721__A1_N _16719_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19611_ _19628_/A VGND VGND VPWR VPWR _19611_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_41_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_83_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16823_ _16823_/A VGND VGND VPWR VPWR _16823_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20250__B2 _20232_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19542_ _19541_/Y _19539_/X _19404_/X _19539_/X VGND VGND VPWR VPWR _19542_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13966_ _13886_/X _13966_/B VGND VGND VPWR VPWR _13966_/X sky130_fd_sc_hd__and2_4
X_16754_ _16752_/Y _16749_/X _16405_/X _16753_/X VGND VGND VPWR VPWR _16754_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_24_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16206__B1 _15949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12917_ _12764_/Y _12917_/B VGND VGND VPWR VPWR _12918_/C sky130_fd_sc_hd__nand2_4
X_15705_ _15713_/A VGND VGND VPWR VPWR _15705_/X sky130_fd_sc_hd__buf_2
XFILLER_62_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16685_ _24480_/Q VGND VGND VPWR VPWR _16685_/Y sky130_fd_sc_hd__inv_2
X_19473_ _23715_/Q VGND VGND VPWR VPWR _22226_/B sky130_fd_sc_hd__inv_2
X_13897_ _13927_/D VGND VGND VPWR VPWR _13897_/X sky130_fd_sc_hd__buf_2
XFILLER_111_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18424_ _24162_/Q VGND VGND VPWR VPWR _18540_/A sky130_fd_sc_hd__inv_2
X_12848_ _25376_/Q VGND VGND VPWR VPWR _12849_/C sky130_fd_sc_hd__inv_2
X_15636_ _21280_/A VGND VGND VPWR VPWR _15636_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15567_ _24908_/Q VGND VGND VPWR VPWR _15567_/Y sky130_fd_sc_hd__inv_2
X_18355_ _18355_/A VGND VGND VPWR VPWR _18355_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12779_ _22895_/A VGND VGND VPWR VPWR _12779_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12243__B2 _24748_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _14502_/X _14516_/X _14474_/A _14517_/X VGND VGND VPWR VPWR _25096_/D sky130_fd_sc_hd__o22a_4
X_17306_ _17344_/A VGND VGND VPWR VPWR _17306_/X sky130_fd_sc_hd__buf_2
XANTENNA__24756__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15498_ _11727_/A VGND VGND VPWR VPWR _15498_/Y sky130_fd_sc_hd__inv_2
X_18286_ _17709_/Y _17702_/A VGND VGND VPWR VPWR _18287_/A sky130_fd_sc_hd__or2_4
X_14449_ _14169_/Y _14448_/X _14395_/X _14448_/X VGND VGND VPWR VPWR _25119_/D sky130_fd_sc_hd__a2bb2o_4
X_17237_ _17237_/A VGND VGND VPWR VPWR _17257_/A sky130_fd_sc_hd__inv_2
XANTENNA__17558__A _17557_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17168_ _17168_/A VGND VGND VPWR VPWR _17169_/A sky130_fd_sc_hd__inv_2
XANTENNA__22463__C1 _22462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16119_ _16117_/Y _16113_/X _15959_/X _16118_/X VGND VGND VPWR VPWR _16119_/X sky130_fd_sc_hd__a2bb2o_4
X_17099_ _17099_/A VGND VGND VPWR VPWR _17099_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16693__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19809_ _19807_/Y _19803_/X _19758_/X _19808_/X VGND VGND VPWR VPWR _19809_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22820_ _22714_/A VGND VGND VPWR VPWR _22820_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_218_0_HCLK clkbuf_8_219_0_HCLK/A VGND VGND VPWR VPWR _24049_/CLK sky130_fd_sc_hd__clkbuf_1
X_22751_ _21422_/X _22746_/X _21826_/X _22750_/Y VGND VGND VPWR VPWR _22751_/X sky130_fd_sc_hd__a211o_4
X_21702_ _21700_/X _21701_/X _21532_/X _24706_/Q _21533_/X VGND VGND VPWR VPWR _21702_/X
+ sky130_fd_sc_hd__a32o_4
X_25470_ _25305_/CLK _12082_/X HRESETn VGND VGND VPWR VPWR _12081_/A sky130_fd_sc_hd__dfrtp_4
X_22682_ _20738_/Y _23126_/A _15602_/Y _22271_/X VGND VGND VPWR VPWR _22682_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24421_ _24427_/CLK _16818_/X HRESETn VGND VGND VPWR VPWR _14969_/A sky130_fd_sc_hd__dfrtp_4
X_21633_ _21633_/A _21625_/X _21632_/X VGND VGND VPWR VPWR _21633_/X sky130_fd_sc_hd__or3_4
XANTENNA__19698__B1 _19553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24497__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24352_ _24356_/CLK _17299_/Y HRESETn VGND VGND VPWR VPWR _23072_/A sky130_fd_sc_hd__dfrtp_4
X_21564_ _18383_/Y _21562_/X _12118_/Y _21561_/X VGND VGND VPWR VPWR _21564_/X sky130_fd_sc_hd__o22a_4
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22374__A _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24426__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23303_ _23271_/A _23303_/B VGND VGND VPWR VPWR _23313_/B sky130_fd_sc_hd__and2_4
X_20515_ _14249_/A _20515_/B _20469_/X _20515_/D VGND VGND VPWR VPWR _20515_/X sky130_fd_sc_hd__or4_4
XFILLER_138_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24283_ _24278_/CLK _17685_/X HRESETn VGND VGND VPWR VPWR _24283_/Q sky130_fd_sc_hd__dfrtp_4
X_21495_ _21994_/A VGND VGND VPWR VPWR _21495_/X sky130_fd_sc_hd__buf_2
XANTENNA__20606__B _17404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23234_ _24530_/Q _22467_/X _22834_/X _23233_/X VGND VGND VPWR VPWR _23235_/C sky130_fd_sc_hd__a211o_4
X_20446_ _20453_/A _20446_/B VGND VGND VPWR VPWR _20446_/X sky130_fd_sc_hd__or2_4
XFILLER_118_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23165_ _23165_/A _23057_/X VGND VGND VPWR VPWR _23169_/B sky130_fd_sc_hd__or2_4
X_20377_ _20377_/A VGND VGND VPWR VPWR _21163_/B sky130_fd_sc_hd__inv_2
XFILLER_134_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16684__B1 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22116_ _14205_/Y _21843_/X _23956_/Q _21351_/B VGND VGND VPWR VPWR _22116_/X sky130_fd_sc_hd__a2bb2o_4
X_23096_ _24760_/Q _23140_/B VGND VGND VPWR VPWR _23096_/X sky130_fd_sc_hd__or2_4
XFILLER_47_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18299__A _18298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22047_ _19543_/Y _21995_/Y _22384_/A _22046_/X VGND VGND VPWR VPWR _22048_/A sky130_fd_sc_hd__a211o_4
XANTENNA__15716__A _15740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18825__A1_N _16501_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14620__A _14620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25285__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_28_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_28_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13820_ _13820_/A VGND VGND VPWR VPWR _13821_/A sky130_fd_sc_hd__buf_2
XANTENNA__13236__A _13227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21980__B2 _21979_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23998_ _24883_/CLK _20685_/Y HRESETn VGND VGND VPWR VPWR _13122_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_21_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23182__B1 _12527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13751_ _13751_/A _13746_/A VGND VGND VPWR VPWR _13752_/A sky130_fd_sc_hd__or2_4
XFILLER_99_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22949_ _15147_/A _22832_/B VGND VGND VPWR VPWR _22952_/B sky130_fd_sc_hd__or2_4
X_12702_ _12731_/A _12729_/A _12728_/A _12735_/A VGND VGND VPWR VPWR _12702_/X sky130_fd_sc_hd__or4_4
XFILLER_44_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16470_ _16469_/Y _16467_/X _16384_/X _16467_/X VGND VGND VPWR VPWR _24562_/D sky130_fd_sc_hd__a2bb2o_4
X_13682_ _13729_/A _13729_/B VGND VGND VPWR VPWR _13683_/B sky130_fd_sc_hd__or2_4
XFILLER_71_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15421_ _15421_/A VGND VGND VPWR VPWR _15421_/Y sky130_fd_sc_hd__inv_2
X_12633_ _12622_/A _12645_/A _12693_/A _12642_/B VGND VGND VPWR VPWR _12636_/B sky130_fd_sc_hd__or4_4
XANTENNA__12225__A1 _25422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24619_ _24345_/CLK _24619_/D HRESETn VGND VGND VPWR VPWR _22940_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_58_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19477__A2_N _19471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15352_ _15298_/C _15352_/B VGND VGND VPWR VPWR _15352_/X sky130_fd_sc_hd__or2_4
X_18140_ _18204_/A _18140_/B VGND VGND VPWR VPWR _18140_/X sky130_fd_sc_hd__or2_4
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12564_ _25389_/Q _12562_/Y _12560_/A _12563_/Y VGND VGND VPWR VPWR _12564_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24914__D _24914_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ _14291_/C _14291_/D _13640_/X _14302_/X VGND VGND VPWR VPWR _14303_/X sky130_fd_sc_hd__a211o_4
XFILLER_12_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18481__B _18481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18071_ _18168_/A _18071_/B VGND VGND VPWR VPWR _18071_/X sky130_fd_sc_hd__or2_4
XANTENNA__24167__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15283_ _15283_/A _15248_/B VGND VGND VPWR VPWR _15283_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15175__B1 _15174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12495_ _12503_/A _12491_/B _12494_/X VGND VGND VPWR VPWR _25425_/D sky130_fd_sc_hd__and3_4
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17022_ _17022_/A VGND VGND VPWR VPWR _17022_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14234_ _14233_/Y _14229_/X _13800_/X _14229_/X VGND VGND VPWR VPWR _14234_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14165_ _14098_/A _14173_/A _25197_/Q _14181_/B VGND VGND VPWR VPWR _14165_/X sky130_fd_sc_hd__or4_4
XFILLER_125_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22460__A2 _21587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12315__A _24826_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13116_ _12311_/Y _13017_/D _13010_/A _13114_/B VGND VGND VPWR VPWR _13116_/X sky130_fd_sc_hd__a211o_4
XFILLER_98_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14096_ scl_oen_o_S4 _20978_/B _14096_/C VGND VGND VPWR VPWR _14096_/X sky130_fd_sc_hd__and3_4
X_18973_ _18971_/Y _18972_/X _17424_/X _18972_/X VGND VGND VPWR VPWR _23890_/D sky130_fd_sc_hd__a2bb2o_4
X_13047_ _25343_/Q _13047_/B VGND VGND VPWR VPWR _13047_/X sky130_fd_sc_hd__or2_4
X_17924_ _17923_/X VGND VGND VPWR VPWR _17924_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15626__A _15561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18002__A _18221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16427__B1 _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17419__A1_N _20662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17855_ _17874_/A _17855_/B _17855_/C VGND VGND VPWR VPWR _24256_/D sky130_fd_sc_hd__and3_4
XFILLER_94_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18937__A _18937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16806_ _24427_/Q VGND VGND VPWR VPWR _16806_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16045__A1_N _16044_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17841__A _17759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17786_ _17786_/A _17786_/B VGND VGND VPWR VPWR _17787_/C sky130_fd_sc_hd__or2_4
X_14998_ _14908_/X _16792_/A _14908_/X _16792_/A VGND VGND VPWR VPWR _15002_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23173__B1 _23172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22459__A _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19525_ _23696_/Q VGND VGND VPWR VPWR _21808_/B sky130_fd_sc_hd__inv_2
XFILLER_130_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16737_ _16736_/Y _16734_/X _16384_/X _16734_/X VGND VGND VPWR VPWR _24461_/D sky130_fd_sc_hd__a2bb2o_4
X_13949_ _13952_/A _13932_/Y _13924_/X _13948_/Y VGND VGND VPWR VPWR _13949_/X sky130_fd_sc_hd__and4_4
Xclkbuf_8_191_0_HCLK clkbuf_7_95_0_HCLK/X VGND VGND VPWR VPWR _25449_/CLK sky130_fd_sc_hd__clkbuf_1
X_19456_ _18110_/B VGND VGND VPWR VPWR _19456_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24937__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16668_ _24487_/Q VGND VGND VPWR VPWR _22984_/A sky130_fd_sc_hd__inv_2
XANTENNA__22490__A1_N _12220_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18407_ _24153_/Q VGND VGND VPWR VPWR _18469_/B sky130_fd_sc_hd__inv_2
XFILLER_37_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_48_0_HCLK clkbuf_8_49_0_HCLK/A VGND VGND VPWR VPWR _25246_/CLK sky130_fd_sc_hd__clkbuf_1
X_15619_ _24887_/Q VGND VGND VPWR VPWR _22407_/A sky130_fd_sc_hd__inv_2
X_19387_ _19386_/Y _19384_/X _19364_/X _19384_/X VGND VGND VPWR VPWR _23745_/D sky130_fd_sc_hd__a2bb2o_4
X_16599_ _24511_/Q VGND VGND VPWR VPWR _16599_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24590__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18338_ _21504_/A _17451_/Y _17476_/A VGND VGND VPWR VPWR _18338_/X sky130_fd_sc_hd__o21a_4
XFILLER_124_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18269_ _13795_/D _18253_/X _16270_/X _23342_/A _18262_/A VGND VGND VPWR VPWR _18269_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14705__A _14705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20300_ _22347_/B _20299_/X _19975_/X _20299_/X VGND VGND VPWR VPWR _23419_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21280_ _21280_/A _21280_/B VGND VGND VPWR VPWR _21286_/B sky130_fd_sc_hd__or2_4
XANTENNA__22922__A _22922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20231_ _17465_/X _18334_/X _20231_/C _19683_/B VGND VGND VPWR VPWR _20232_/A sky130_fd_sc_hd__or4_4
X_20162_ _21616_/B _20161_/X _20096_/X _20161_/X VGND VGND VPWR VPWR _23471_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20093_ _20091_/Y _20086_/X _20092_/X _20086_/X VGND VGND VPWR VPWR _23496_/D sky130_fd_sc_hd__a2bb2o_4
X_24970_ _24980_/CLK _24970_/D HRESETn VGND VGND VPWR VPWR _24970_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23921_ _23959_/CLK _23921_/D HRESETn VGND VGND VPWR VPWR _23921_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14968__A2_N _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23852_ _24398_/CLK _19087_/X VGND VGND VPWR VPWR _19083_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_66_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22803_ _24550_/Q _22421_/X _22526_/X VGND VGND VPWR VPWR _22803_/X sky130_fd_sc_hd__o21a_4
XFILLER_26_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23783_ _23846_/CLK _23783_/D VGND VGND VPWR VPWR _23783_/Q sky130_fd_sc_hd__dfxtp_4
X_20995_ _20996_/A _20995_/B _23968_/Q VGND VGND VPWR VPWR _20995_/X sky130_fd_sc_hd__and3_4
XFILLER_111_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25522_ _24275_/CLK _25522_/D HRESETn VGND VGND VPWR VPWR _25522_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24678__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22734_ _16501_/A _22525_/X _22527_/X VGND VGND VPWR VPWR _22734_/X sky130_fd_sc_hd__o21a_4
XFILLER_111_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24607__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25453_ _24383_/CLK _25453_/D HRESETn VGND VGND VPWR VPWR _25453_/Q sky130_fd_sc_hd__dfrtp_4
X_22665_ _16832_/Y _21413_/X _21573_/X _22664_/X VGND VGND VPWR VPWR _22665_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22816__B _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24404_ _24435_/CLK _24404_/D HRESETn VGND VGND VPWR VPWR _16850_/A sky130_fd_sc_hd__dfrtp_4
X_21616_ _21616_/A _21616_/B VGND VGND VPWR VPWR _21619_/B sky130_fd_sc_hd__or2_4
X_25384_ _25385_/CLK _12873_/X HRESETn VGND VGND VPWR VPWR _12871_/A sky130_fd_sc_hd__dfrtp_4
X_22596_ _22544_/X _22595_/X _22125_/X _25518_/Q _22922_/A VGND VGND VPWR VPWR _22596_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__11966__B1 _11965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24260__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24335_ _24334_/CLK _24335_/D HRESETn VGND VGND VPWR VPWR _24335_/Q sky130_fd_sc_hd__dfrtp_4
X_21547_ _21547_/A VGND VGND VPWR VPWR _21547_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20150__B1 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12280_ _12280_/A VGND VGND VPWR VPWR _12280_/Y sky130_fd_sc_hd__inv_2
X_24266_ _24692_/CLK _17815_/X HRESETn VGND VGND VPWR VPWR _16900_/A sky130_fd_sc_hd__dfrtp_4
X_21478_ _21478_/A VGND VGND VPWR VPWR _21484_/A sky130_fd_sc_hd__buf_2
XFILLER_4_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23217_ _23106_/X _23216_/X _23040_/X _24731_/Q _21520_/X VGND VGND VPWR VPWR _23217_/X
+ sky130_fd_sc_hd__a32o_4
X_20429_ _20428_/X VGND VGND VPWR VPWR _20429_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24197_ _24197_/CLK _18330_/Y HRESETn VGND VGND VPWR VPWR _24197_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25466__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21448__A _21455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23148_ _23106_/X _23147_/X _23040_/X _24729_/Q _22972_/X VGND VGND VPWR VPWR _23148_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20352__A _20339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15970_ _15966_/X _15969_/X _11800_/A _24750_/Q _15967_/X VGND VGND VPWR VPWR _24750_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_27_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23079_ _16660_/Y _22824_/X _15577_/Y _22827_/X VGND VGND VPWR VPWR _23079_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16409__B1 _16408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14921_ _25002_/Q VGND VGND VPWR VPWR _15064_/A sky130_fd_sc_hd__inv_2
XFILLER_49_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15165__B _15165_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17640_ _17525_/Y _17639_/X VGND VGND VPWR VPWR _17641_/B sky130_fd_sc_hd__or2_4
XANTENNA__17661__A _17557_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14852_ _25035_/Q _14814_/X _25035_/Q _14814_/X VGND VGND VPWR VPWR _14852_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13803_ _15986_/A VGND VGND VPWR VPWR _13803_/X sky130_fd_sc_hd__buf_2
X_14783_ _14783_/A VGND VGND VPWR VPWR _14783_/Y sky130_fd_sc_hd__inv_2
X_17571_ _17571_/A VGND VGND VPWR VPWR _17571_/Y sky130_fd_sc_hd__inv_2
X_11995_ _11994_/X VGND VGND VPWR VPWR _11995_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21705__B2 _23100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19310_ _19038_/A _19014_/B _19399_/C VGND VGND VPWR VPWR _19310_/X sky130_fd_sc_hd__or3_4
Xclkbuf_8_201_0_HCLK clkbuf_8_201_0_HCLK/A VGND VGND VPWR VPWR _24806_/CLK sky130_fd_sc_hd__clkbuf_1
X_13734_ _25267_/Q VGND VGND VPWR VPWR _13735_/A sky130_fd_sc_hd__inv_2
X_16522_ _16520_/Y _16516_/X _16521_/X _16516_/X VGND VGND VPWR VPWR _24541_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_7_0_HCLK clkbuf_8_7_0_HCLK/A VGND VGND VPWR VPWR _23478_/CLK sky130_fd_sc_hd__clkbuf_1
X_19241_ _23796_/Q VGND VGND VPWR VPWR _22354_/B sky130_fd_sc_hd__inv_2
XFILLER_95_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24348__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13665_ _13664_/X VGND VGND VPWR VPWR _20922_/B sky130_fd_sc_hd__buf_2
X_16453_ _16453_/A _16453_/B _15533_/Y _11732_/A VGND VGND VPWR VPWR _16454_/A sky130_fd_sc_hd__or4_4
XANTENNA__15396__B1 _15339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12616_ _12704_/A _12616_/B _12728_/A _12529_/Y VGND VGND VPWR VPWR _12616_/X sky130_fd_sc_hd__or4_4
X_15404_ _15392_/A _15408_/A VGND VGND VPWR VPWR _15404_/Y sky130_fd_sc_hd__nand2_4
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16384_ HWDATA[28] VGND VGND VPWR VPWR _16384_/X sky130_fd_sc_hd__buf_2
X_19172_ _19171_/Y _19167_/X _19149_/X _19153_/Y VGND VGND VPWR VPWR _19172_/X sky130_fd_sc_hd__a2bb2o_4
X_13596_ _12095_/A _16453_/A _13813_/A _13777_/A VGND VGND VPWR VPWR _14433_/A sky130_fd_sc_hd__or4_4
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15335_ _15334_/X VGND VGND VPWR VPWR _24989_/D sky130_fd_sc_hd__inv_2
X_18123_ _18187_/A _18123_/B VGND VGND VPWR VPWR _18124_/C sky130_fd_sc_hd__or2_4
X_12547_ _25417_/Q _24871_/Q _12636_/A _12546_/Y VGND VGND VPWR VPWR _12557_/A sky130_fd_sc_hd__o22a_4
XANTENNA__20141__B1 _20096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15266_ _14942_/Y _15272_/A VGND VGND VPWR VPWR _15267_/B sky130_fd_sc_hd__or2_4
X_18054_ _18088_/A VGND VGND VPWR VPWR _18054_/X sky130_fd_sc_hd__buf_2
X_12478_ _12282_/C _12477_/X _12412_/A _12474_/B VGND VGND VPWR VPWR _12479_/A sky130_fd_sc_hd__a211o_4
X_14217_ _14216_/Y _14201_/A _13800_/X _14201_/A VGND VGND VPWR VPWR _14217_/X sky130_fd_sc_hd__a2bb2o_4
X_17005_ _24388_/Q VGND VGND VPWR VPWR _17005_/Y sky130_fd_sc_hd__inv_2
X_15197_ _15197_/A _15194_/X VGND VGND VPWR VPWR _15198_/C sky130_fd_sc_hd__or2_4
XANTENNA__19834__B1 _19790_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23983__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14148_ _14147_/X VGND VGND VPWR VPWR _14148_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25136__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14079_ _13990_/C _14065_/X _14078_/X _13998_/X _14076_/X VGND VGND VPWR VPWR _14079_/X
+ sky130_fd_sc_hd__a32o_4
X_18956_ _18954_/Y _18952_/X _18955_/X _18952_/X VGND VGND VPWR VPWR _18956_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17907_ _17909_/A _17894_/X VGND VGND VPWR VPWR _17907_/X sky130_fd_sc_hd__or2_4
XFILLER_117_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18887_ _18869_/X _18883_/X _24110_/Q _20974_/A _18886_/X VGND VGND VPWR VPWR _24111_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13882__B1 _23428_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17838_ _17753_/Y _17837_/X VGND VGND VPWR VPWR _17841_/B sky130_fd_sc_hd__or2_4
Xclkbuf_6_11_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_94_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16820__B1 HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17769_ _17738_/X _17767_/X _17768_/Y VGND VGND VPWR VPWR _24276_/D sky130_fd_sc_hd__and3_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19508_ _19506_/Y _19507_/X _11952_/X _19507_/X VGND VGND VPWR VPWR _19508_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13604__A _14645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24771__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20780_ _20779_/Y _20776_/Y _20783_/B VGND VGND VPWR VPWR _20780_/X sky130_fd_sc_hd__o21a_4
XFILLER_62_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21821__A _21821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24089__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24700__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19439_ _19437_/Y _19438_/X _19370_/X _19438_/X VGND VGND VPWR VPWR _19439_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24018__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22450_ _18230_/A VGND VGND VPWR VPWR _22613_/B sky130_fd_sc_hd__buf_2
X_21401_ _21391_/A _21399_/X _21400_/X VGND VGND VPWR VPWR _21401_/X sky130_fd_sc_hd__and3_4
X_22381_ _21507_/Y _22352_/X _13775_/X _22380_/X VGND VGND VPWR VPWR _22381_/Y sky130_fd_sc_hd__a22oi_4
X_24120_ _24120_/CLK _18805_/X HRESETn VGND VGND VPWR VPWR _18623_/A sky130_fd_sc_hd__dfrtp_4
X_21332_ _21331_/X VGND VGND VPWR VPWR _21332_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24051_ _24487_/CLK _20917_/X HRESETn VGND VGND VPWR VPWR _24051_/Q sky130_fd_sc_hd__dfrtp_4
X_21263_ _23669_/Q _20318_/X _23685_/Q _21200_/B VGND VGND VPWR VPWR _21263_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19825__B1 _19777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23002_ _23002_/A _22990_/Y _23002_/C _23002_/D VGND VGND VPWR VPWR _23002_/X sky130_fd_sc_hd__or4_4
X_20214_ _23451_/Q VGND VGND VPWR VPWR _20214_/Y sky130_fd_sc_hd__inv_2
X_21194_ _21194_/A _21194_/B _21194_/C VGND VGND VPWR VPWR _21194_/X sky130_fd_sc_hd__and3_4
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20145_ _20144_/Y _20140_/X _20123_/X _20140_/A VGND VGND VPWR VPWR _20145_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24953_ _24950_/CLK _15451_/X HRESETn VGND VGND VPWR VPWR _13909_/A sky130_fd_sc_hd__dfrtp_4
X_20076_ _20076_/A VGND VGND VPWR VPWR _22371_/B sky130_fd_sc_hd__inv_2
XANTENNA__20900__A _20900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18800__A1 _18792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24859__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23904_ _23904_/CLK _18935_/X VGND VGND VPWR VPWR _13347_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21715__B _21549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24884_ _24885_/CLK _24884_/D HRESETn VGND VGND VPWR VPWR _15629_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23835_ _23884_/CLK _23835_/D VGND VGND VPWR VPWR _19132_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_26_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16505__A1_N _16503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25289__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11780_ _25527_/Q VGND VGND VPWR VPWR _11780_/Y sky130_fd_sc_hd__inv_2
X_23766_ _23660_/CLK _23766_/D VGND VGND VPWR VPWR _23766_/Q sky130_fd_sc_hd__dfxtp_4
X_20978_ _20978_/A _20978_/B _20977_/C VGND VGND VPWR VPWR _20979_/A sky130_fd_sc_hd__or3_4
XFILLER_82_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21731__A _22524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24441__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25505_ _25503_/CLK _25505_/D HRESETn VGND VGND VPWR VPWR _25505_/Q sky130_fd_sc_hd__dfrtp_4
X_22717_ _22425_/X _22713_/X _22714_/X _22716_/Y VGND VGND VPWR VPWR _22718_/B sky130_fd_sc_hd__o22a_4
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23697_ _24926_/CLK _19524_/X VGND VGND VPWR VPWR _19523_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13450_ _13450_/A _13448_/X _13450_/C VGND VGND VPWR VPWR _13454_/B sky130_fd_sc_hd__and3_4
XFILLER_16_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18743__C _18743_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_31_0_HCLK clkbuf_8_31_0_HCLK/A VGND VGND VPWR VPWR _24364_/CLK sky130_fd_sc_hd__clkbuf_1
X_25436_ _25436_/CLK _12451_/Y HRESETn VGND VGND VPWR VPWR _12187_/A sky130_fd_sc_hd__dfrtp_4
X_22648_ _15709_/A _22647_/X _22130_/C _24820_/Q _22677_/B VGND VGND VPWR VPWR _22649_/B
+ sky130_fd_sc_hd__a32o_4
X_12401_ _12389_/A _12401_/B _12400_/X VGND VGND VPWR VPWR _12401_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_94_0_HCLK clkbuf_8_95_0_HCLK/A VGND VGND VPWR VPWR _24120_/CLK sky130_fd_sc_hd__clkbuf_1
X_13381_ _13413_/A _13379_/X _13381_/C VGND VGND VPWR VPWR _13382_/C sky130_fd_sc_hd__and3_4
XFILLER_90_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25367_ _25356_/CLK _12938_/Y HRESETn VGND VGND VPWR VPWR _25367_/Q sky130_fd_sc_hd__dfrtp_4
X_22579_ _20867_/Y _21588_/X _20728_/Y _22988_/A VGND VGND VPWR VPWR _22579_/X sky130_fd_sc_hd__o22a_4
X_15120_ _15120_/A _15113_/X _15116_/X _15120_/D VGND VGND VPWR VPWR _15120_/X sky130_fd_sc_hd__or4_4
X_12332_ _12330_/A _24816_/Q _13092_/A _12331_/Y VGND VGND VPWR VPWR _12332_/X sky130_fd_sc_hd__o22a_4
X_24318_ _24318_/CLK _17426_/X HRESETn VGND VGND VPWR VPWR _17423_/A sky130_fd_sc_hd__dfrtp_4
X_25298_ _25301_/CLK _25298_/D HRESETn VGND VGND VPWR VPWR _25298_/Q sky130_fd_sc_hd__dfrtp_4
X_15051_ _24459_/Q VGND VGND VPWR VPWR _15051_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12263_ _12263_/A VGND VGND VPWR VPWR _12263_/Y sky130_fd_sc_hd__inv_2
X_24249_ _24673_/CLK _17876_/Y HRESETn VGND VGND VPWR VPWR _17745_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22415__A2 _22288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19816__B1 _19721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14002_ _14002_/A _13983_/A _25220_/Q _25219_/Q VGND VGND VPWR VPWR _14002_/X sky130_fd_sc_hd__or4_4
XANTENNA__22281__B _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12194_ _23178_/A VGND VGND VPWR VPWR _12194_/Y sky130_fd_sc_hd__inv_2
X_18810_ _18799_/A _18803_/B _18810_/C VGND VGND VPWR VPWR _24118_/D sky130_fd_sc_hd__and3_4
X_19790_ _19790_/A VGND VGND VPWR VPWR _19790_/X sky130_fd_sc_hd__buf_2
X_18741_ _18740_/X VGND VGND VPWR VPWR _24135_/D sky130_fd_sc_hd__inv_2
X_15953_ _12259_/Y _15945_/X _15952_/X _15945_/X VGND VGND VPWR VPWR _24757_/D sky130_fd_sc_hd__a2bb2o_4
X_14904_ _24422_/Q VGND VGND VPWR VPWR _14904_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18672_ _24139_/Q VGND VGND VPWR VPWR _18672_/Y sky130_fd_sc_hd__inv_2
X_15884_ _12765_/Y _15882_/X _11788_/X _15882_/X VGND VGND VPWR VPWR _15884_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17623_ _17623_/A VGND VGND VPWR VPWR _17623_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24529__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14835_ _14809_/A VGND VGND VPWR VPWR _14835_/X sky130_fd_sc_hd__buf_2
XFILLER_40_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17554_ _17837_/A VGND VGND VPWR VPWR _17624_/A sky130_fd_sc_hd__buf_2
X_11978_ _11976_/X VGND VGND VPWR VPWR _11978_/Y sky130_fd_sc_hd__inv_2
X_14766_ _13743_/A _13742_/A VGND VGND VPWR VPWR _14766_/X sky130_fd_sc_hd__and2_4
XANTENNA__22351__A1 _17722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22737__A _24787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16505_ _16503_/Y _16499_/X _16231_/X _16504_/X VGND VGND VPWR VPWR _24548_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24182__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13717_ _13689_/B _13707_/X _13716_/Y _13714_/X _11685_/A VGND VGND VPWR VPWR _25276_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_60_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14697_ _14697_/A _14697_/B VGND VGND VPWR VPWR _14698_/D sky130_fd_sc_hd__and2_4
X_17485_ _17457_/A _17483_/X _17457_/Y _17484_/Y VGND VGND VPWR VPWR _17485_/X sky130_fd_sc_hd__o22a_4
X_19224_ _13211_/B VGND VGND VPWR VPWR _19224_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16436_ _24571_/Q VGND VGND VPWR VPWR _16436_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13648_ _24056_/Q _20931_/A VGND VGND VPWR VPWR _13648_/X sky130_fd_sc_hd__or2_4
XFILLER_73_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11879__A _11700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19155_ _19017_/X VGND VGND VPWR VPWR _19155_/X sky130_fd_sc_hd__buf_2
XANTENNA__20114__B1 _20089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13579_ _25079_/Q VGND VGND VPWR VPWR _14592_/A sky130_fd_sc_hd__inv_2
X_16367_ _16365_/Y _16282_/A _16366_/X _16282_/A VGND VGND VPWR VPWR _16367_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14255__A _14255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_2_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18106_ _18217_/A _18102_/X _18106_/C VGND VGND VPWR VPWR _18114_/B sky130_fd_sc_hd__or3_4
XANTENNA__25388__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15318_ _15318_/A _15312_/B _15317_/X VGND VGND VPWR VPWR _15318_/X sky130_fd_sc_hd__or3_4
X_16298_ _16295_/Y _16296_/X _16297_/X _16296_/X VGND VGND VPWR VPWR _24625_/D sky130_fd_sc_hd__a2bb2o_4
X_19086_ _19098_/A VGND VGND VPWR VPWR _19086_/X sky130_fd_sc_hd__buf_2
XANTENNA__25317__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18037_ _18180_/A _23890_/Q VGND VGND VPWR VPWR _18038_/C sky130_fd_sc_hd__or2_4
X_15249_ _15249_/A _15249_/B VGND VGND VPWR VPWR _15272_/A sky130_fd_sc_hd__or2_4
XANTENNA__15541__B1 HADDR[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21090__B2 _21729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19988_ _11941_/A VGND VGND VPWR VPWR _19988_/X sky130_fd_sc_hd__buf_2
XFILLER_45_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18939_ _13411_/B VGND VGND VPWR VPWR _18939_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21816__A _24198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21950_ _21950_/A VGND VGND VPWR VPWR _21950_/X sky130_fd_sc_hd__buf_2
XFILLER_55_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24952__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20901_ _20901_/A VGND VGND VPWR VPWR _20901_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21881_ _21886_/A _21881_/B VGND VGND VPWR VPWR _21881_/X sky130_fd_sc_hd__or2_4
XFILLER_55_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18609__A1_N _16597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23620_ _23635_/CLK _23620_/D VGND VGND VPWR VPWR _13170_/B sky130_fd_sc_hd__dfxtp_4
X_20832_ _13657_/B VGND VGND VPWR VPWR _20832_/Y sky130_fd_sc_hd__inv_2
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21145__A2 _14220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22647__A _24748_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23551_ _25433_/CLK _19944_/X VGND VGND VPWR VPWR _19942_/A sky130_fd_sc_hd__dfxtp_4
X_20763_ _13119_/D _20758_/X _20767_/B VGND VGND VPWR VPWR _20763_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16645__A _16645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22502_ _20717_/Y _22988_/A _20856_/Y _22790_/A VGND VGND VPWR VPWR _22502_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_18_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23482_ _23498_/CLK _20134_/X VGND VGND VPWR VPWR _20132_/A sky130_fd_sc_hd__dfxtp_4
X_20694_ _13127_/B VGND VGND VPWR VPWR _20694_/Y sky130_fd_sc_hd__inv_2
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25221_ _25043_/CLK _14082_/X HRESETn VGND VGND VPWR VPWR _25221_/Q sky130_fd_sc_hd__dfrtp_4
X_22433_ _22433_/A VGND VGND VPWR VPWR _22434_/D sky130_fd_sc_hd__inv_2
XANTENNA__21853__B1 _21103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25152_ _24109_/CLK _14342_/X HRESETn VGND VGND VPWR VPWR _25152_/Q sky130_fd_sc_hd__dfrtp_4
X_22364_ _22068_/A _22364_/B VGND VGND VPWR VPWR _22364_/X sky130_fd_sc_hd__or2_4
XANTENNA__22382__A _21821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25058__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24103_ _24109_/CLK MSI_S3 HRESETn VGND VGND VPWR VPWR _24103_/Q sky130_fd_sc_hd__dfrtp_4
X_21315_ _21314_/X VGND VGND VPWR VPWR _21316_/A sky130_fd_sc_hd__buf_2
XANTENNA__15532__B1 HADDR[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25083_ _24376_/CLK _14583_/X HRESETn VGND VGND VPWR VPWR _13570_/A sky130_fd_sc_hd__dfrtp_4
X_22295_ _24541_/Q _22590_/B _22885_/A VGND VGND VPWR VPWR _22295_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16380__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24034_ _24649_/CLK _20840_/Y HRESETn VGND VGND VPWR VPWR _24034_/Q sky130_fd_sc_hd__dfrtp_4
X_21246_ _21249_/A _19927_/Y VGND VGND VPWR VPWR _21247_/C sky130_fd_sc_hd__or2_4
XANTENNA__23070__A2 _22393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21177_ _21185_/A _21177_/B VGND VGND VPWR VPWR _21178_/C sky130_fd_sc_hd__or2_4
XFILLER_63_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20128_ _20140_/A VGND VGND VPWR VPWR _20128_/X sky130_fd_sc_hd__buf_2
X_12950_ _12944_/C _12949_/X _12884_/A _12945_/Y VGND VGND VPWR VPWR _12951_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24693__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20059_ _23510_/Q VGND VGND VPWR VPWR _20059_/Y sky130_fd_sc_hd__inv_2
X_24936_ _25508_/CLK _24936_/D HRESETn VGND VGND VPWR VPWR _24936_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11901_ _11901_/A VGND VGND VPWR VPWR _11902_/B sky130_fd_sc_hd__buf_2
XFILLER_100_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24622__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12881_ _12881_/A _12879_/X _12881_/C VGND VGND VPWR VPWR _25382_/D sky130_fd_sc_hd__and3_4
XFILLER_34_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24867_ _24865_/CLK _15726_/X HRESETn VGND VGND VPWR VPWR _24867_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11832_ HWDATA[7] VGND VGND VPWR VPWR _13835_/A sky130_fd_sc_hd__buf_2
X_14620_ _14620_/A _14620_/B _13598_/X _14620_/D VGND VGND VPWR VPWR _14620_/X sky130_fd_sc_hd__and4_4
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23818_ _23818_/CLK _23818_/D VGND VGND VPWR VPWR _19180_/A sky130_fd_sc_hd__dfxtp_4
X_24798_ _24830_/CLK _15874_/X HRESETn VGND VGND VPWR VPWR _24798_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22557__A _21582_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ HSEL VGND VGND VPWR VPWR _14551_/X sky130_fd_sc_hd__buf_2
XFILLER_26_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11763_/A VGND VGND VPWR VPWR _11763_/Y sky130_fd_sc_hd__inv_2
XPHY_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23749_ _23446_/CLK _23749_/D VGND VGND VPWR VPWR _18196_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16555__A _24529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _11990_/Y _13498_/X _11833_/X _13501_/X VGND VGND VPWR VPWR _25301_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14480_/Y _14476_/X _14418_/X _14481_/X VGND VGND VPWR VPWR _25106_/D sky130_fd_sc_hd__a2bb2o_4
X_17270_ _17231_/X VGND VGND VPWR VPWR _17279_/A sky130_fd_sc_hd__inv_2
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20895__B2 _20886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _24215_/Q VGND VGND VPWR VPWR _11694_/Y sky130_fd_sc_hd__inv_2
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13433_ _17452_/B _23853_/Q VGND VGND VPWR VPWR _13433_/X sky130_fd_sc_hd__or2_4
X_16221_ _22809_/A VGND VGND VPWR VPWR _16221_/Y sky130_fd_sc_hd__inv_2
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25419_ _25400_/CLK _12627_/X HRESETn VGND VGND VPWR VPWR _25419_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15771__B1 _14470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25481__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16152_ _16125_/X VGND VGND VPWR VPWR _16152_/X sky130_fd_sc_hd__buf_2
X_13364_ _13428_/A _13362_/X _13363_/X VGND VGND VPWR VPWR _13364_/X sky130_fd_sc_hd__and3_4
XANTENNA__25410__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12315_ _24826_/Q VGND VGND VPWR VPWR _12315_/Y sky130_fd_sc_hd__inv_2
X_15103_ _24987_/Q _24591_/Q _15338_/A _15102_/Y VGND VGND VPWR VPWR _15107_/C sky130_fd_sc_hd__o22a_4
X_16083_ _23310_/A VGND VGND VPWR VPWR _16083_/Y sky130_fd_sc_hd__inv_2
X_13295_ _13200_/X _13276_/X _13294_/X _25319_/Q _11965_/X VGND VGND VPWR VPWR _13295_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_127_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15034_ _15193_/A _16745_/A _15193_/A _16745_/A VGND VGND VPWR VPWR _15034_/X sky130_fd_sc_hd__a2bb2o_4
X_19911_ _19923_/A VGND VGND VPWR VPWR _19911_/X sky130_fd_sc_hd__buf_2
X_12246_ _25437_/Q VGND VGND VPWR VPWR _12286_/B sky130_fd_sc_hd__inv_2
X_19842_ _21223_/B _19836_/X _19841_/X _19836_/A VGND VGND VPWR VPWR _23589_/D sky130_fd_sc_hd__a2bb2o_4
X_12177_ _12474_/A VGND VGND VPWR VPWR _12475_/A sky130_fd_sc_hd__inv_2
XFILLER_1_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19773_ _23612_/Q VGND VGND VPWR VPWR _19773_/Y sky130_fd_sc_hd__inv_2
X_16985_ _16985_/A VGND VGND VPWR VPWR _16985_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18724_ _18724_/A _18724_/B _18724_/C VGND VGND VPWR VPWR _18725_/A sky130_fd_sc_hd__or3_4
XFILLER_114_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15936_ _15930_/X _15935_/X HWDATA[30] _24765_/Q _15933_/X VGND VGND VPWR VPWR _15936_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_3_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18010__A _18010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22572__A1 _24444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24363__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18655_ _16613_/Y _24117_/Q _24530_/Q _18654_/Y VGND VGND VPWR VPWR _18655_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15867_ _15863_/A VGND VGND VPWR VPWR _15900_/A sky130_fd_sc_hd__inv_2
XFILLER_92_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17606_ _17600_/C _17604_/A VGND VGND VPWR VPWR _17606_/X sky130_fd_sc_hd__or2_4
X_14818_ _14817_/X VGND VGND VPWR VPWR _14819_/B sky130_fd_sc_hd__inv_2
X_18586_ _18418_/Y _18585_/X VGND VGND VPWR VPWR _18588_/B sky130_fd_sc_hd__or2_4
XFILLER_75_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15798_ _15829_/A VGND VGND VPWR VPWR _15809_/A sky130_fd_sc_hd__buf_2
XANTENNA__14262__B1 _13837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17537_ _17533_/X _17537_/B _17537_/C _17536_/X VGND VGND VPWR VPWR _17551_/B sky130_fd_sc_hd__or4_4
X_14749_ _14749_/A VGND VGND VPWR VPWR _14749_/X sky130_fd_sc_hd__buf_2
XANTENNA__16465__A _24563_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17468_ _24195_/Q _24194_/Q VGND VGND VPWR VPWR _17468_/X sky130_fd_sc_hd__and2_4
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19207_ _19205_/Y _19203_/X _19206_/X _19203_/X VGND VGND VPWR VPWR _23809_/D sky130_fd_sc_hd__a2bb2o_4
X_16419_ _16433_/A VGND VGND VPWR VPWR _16419_/X sky130_fd_sc_hd__buf_2
XANTENNA__15762__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19776__A _19793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17399_ _17399_/A _17399_/B VGND VGND VPWR VPWR _17402_/B sky130_fd_sc_hd__or2_4
XFILLER_125_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19138_ _19135_/Y _19130_/X _19136_/X _19137_/X VGND VGND VPWR VPWR _23834_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17296__A _17239_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19069_ _19067_/Y _19063_/X _18997_/X _19068_/X VGND VGND VPWR VPWR _23858_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15514__B1 HADDR[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21100_ _21064_/X _21065_/X _21082_/X _21094_/X _21099_/X VGND VGND VPWR VPWR _21274_/C
+ sky130_fd_sc_hd__a32o_4
X_22080_ _14693_/A _22075_/X _22076_/X _22077_/X _22079_/X VGND VGND VPWR VPWR _22080_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_114_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21031_ _15649_/A _21074_/B VGND VGND VPWR VPWR _21031_/X sky130_fd_sc_hd__and2_4
XFILLER_102_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13828__B1 _11818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15544__A _21582_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22982_ _17252_/C _22908_/X _25376_/Q _22909_/X VGND VGND VPWR VPWR _22982_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12500__B1 _12394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21933_ _21469_/A _21922_/X _21932_/X VGND VGND VPWR VPWR _21933_/X sky130_fd_sc_hd__or3_4
X_24721_ _24720_/CLK _24721_/D HRESETn VGND VGND VPWR VPWR _16029_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24033__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24652_ _24162_/CLK _16220_/X HRESETn VGND VGND VPWR VPWR _22878_/A sky130_fd_sc_hd__dfrtp_4
X_21864_ _22664_/B VGND VGND VPWR VPWR _23005_/C sky130_fd_sc_hd__buf_2
X_23603_ _23618_/CLK _19806_/X VGND VGND VPWR VPWR _13253_/B sky130_fd_sc_hd__dfxtp_4
X_20815_ _20814_/X VGND VGND VPWR VPWR _20815_/X sky130_fd_sc_hd__buf_2
XFILLER_93_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24583_ _24572_/CLK _16415_/X HRESETn VGND VGND VPWR VPWR _24583_/Q sky130_fd_sc_hd__dfrtp_4
X_21795_ _21456_/A _21795_/B VGND VGND VPWR VPWR _21795_/X sky130_fd_sc_hd__or2_4
XANTENNA__12803__B2 _22708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19192__B1 _19191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23534_ _23711_/CLK _19996_/X VGND VGND VPWR VPWR _23534_/Q sky130_fd_sc_hd__dfxtp_4
X_20746_ _24012_/Q _20740_/X _20745_/Y VGND VGND VPWR VPWR _20746_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25239__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15753__B1 _24853_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23465_ _23581_/CLK _23465_/D VGND VGND VPWR VPWR _23465_/Q sky130_fd_sc_hd__dfxtp_4
X_20677_ _20676_/X VGND VGND VPWR VPWR _20677_/X sky130_fd_sc_hd__buf_2
XANTENNA__25057__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12408__A _12291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25204_ _25205_/CLK _25204_/D HRESETn VGND VGND VPWR VPWR _14115_/A sky130_fd_sc_hd__dfrtp_4
X_22416_ _23281_/A _22409_/Y _22412_/X _22413_/X _22415_/X VGND VGND VPWR VPWR _22417_/D
+ sky130_fd_sc_hd__o32a_4
X_23396_ _23396_/CLK _23396_/D VGND VGND VPWR VPWR _23396_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_104_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_105_0_HCLK clkbuf_7_52_0_HCLK/X VGND VGND VPWR VPWR _24612_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_137_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25135_ _25178_/CLK _25135_/D HRESETn VGND VGND VPWR VPWR _25135_/Q sky130_fd_sc_hd__dfrtp_4
X_22347_ _21458_/A _22347_/B VGND VGND VPWR VPWR _22347_/X sky130_fd_sc_hd__or2_4
XANTENNA__15505__B1 HADDR[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_168_0_HCLK clkbuf_7_84_0_HCLK/X VGND VGND VPWR VPWR _23682_/CLK sky130_fd_sc_hd__clkbuf_1
X_12100_ _13533_/D _13496_/B _12066_/X _12100_/D VGND VGND VPWR VPWR _12101_/A sky130_fd_sc_hd__or4_4
X_13080_ _12993_/A _13107_/A _13106_/A _13113_/A VGND VGND VPWR VPWR _13081_/B sky130_fd_sc_hd__or4_4
X_25066_ _25054_/CLK _14635_/X HRESETn VGND VGND VPWR VPWR _14632_/A sky130_fd_sc_hd__dfrtp_4
X_22278_ _21581_/X VGND VGND VPWR VPWR _22278_/X sky130_fd_sc_hd__buf_2
XANTENNA__22840__A _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21159__C _21158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12031_ _25481_/Q VGND VGND VPWR VPWR _12031_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21054__A1 _24701_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24017_ _24868_/CLK _20769_/X HRESETn VGND VGND VPWR VPWR _13120_/B sky130_fd_sc_hd__dfrtp_4
X_21229_ _21252_/A _21229_/B VGND VGND VPWR VPWR _21229_/X sky130_fd_sc_hd__or2_4
XANTENNA__24874__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24803__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16770_ _16773_/A VGND VGND VPWR VPWR _16770_/X sky130_fd_sc_hd__buf_2
X_13982_ _13982_/A VGND VGND VPWR VPWR _13984_/C sky130_fd_sc_hd__inv_2
XANTENNA__13295__B2 _11965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15721_ _15721_/A VGND VGND VPWR VPWR _15721_/X sky130_fd_sc_hd__buf_2
XFILLER_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12933_ _12933_/A VGND VGND VPWR VPWR _12933_/Y sky130_fd_sc_hd__inv_2
X_24919_ _25433_/CLK _15530_/X HRESETn VGND VGND VPWR VPWR _24919_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18440_ _24165_/Q VGND VGND VPWR VPWR _18524_/A sky130_fd_sc_hd__inv_2
XANTENNA__17430__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15652_ _15662_/A _15662_/B _11732_/A _15652_/D VGND VGND VPWR VPWR _15653_/A sky130_fd_sc_hd__or4_4
X_12864_ _12864_/A _12840_/Y _12863_/X VGND VGND VPWR VPWR _12864_/X sky130_fd_sc_hd__or3_4
XANTENNA__24917__D _15534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14603_ _14564_/X _14601_/Y _14599_/X _14602_/X _13559_/A VGND VGND VPWR VPWR _14603_/X
+ sky130_fd_sc_hd__a32o_4
X_11815_ _25518_/Q VGND VGND VPWR VPWR _11815_/Y sky130_fd_sc_hd__inv_2
X_18371_ _18371_/A VGND VGND VPWR VPWR _18377_/A sky130_fd_sc_hd__inv_2
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12795_ _21414_/A VGND VGND VPWR VPWR _12795_/Y sky130_fd_sc_hd__inv_2
X_15583_ _15583_/A VGND VGND VPWR VPWR _15583_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16285__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17254_/A _17321_/X VGND VGND VPWR VPWR _17322_/Y sky130_fd_sc_hd__nand2_4
XPHY_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ HWDATA[30] VGND VGND VPWR VPWR _11746_/X sky130_fd_sc_hd__buf_2
X_14534_ _20531_/A _14071_/X VGND VGND VPWR VPWR _14534_/X sky130_fd_sc_hd__and2_4
XFILLER_30_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ _24344_/Q VGND VGND VPWR VPWR _17253_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _11677_/A VGND VGND VPWR VPWR _11677_/Y sky130_fd_sc_hd__inv_2
X_14465_ _14465_/A VGND VGND VPWR VPWR _14465_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22609__A2 _22525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15744__B1 _24857_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16204_ _23068_/A VGND VGND VPWR VPWR _16204_/Y sky130_fd_sc_hd__inv_2
X_13416_ _13316_/A _19678_/A VGND VGND VPWR VPWR _13416_/X sky130_fd_sc_hd__or2_4
XFILLER_70_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_64_0_HCLK clkbuf_6_32_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_64_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14396_ _14393_/Y _14394_/X _14395_/X _14384_/X VGND VGND VPWR VPWR _14396_/X sky130_fd_sc_hd__a2bb2o_4
X_17184_ _17184_/A VGND VGND VPWR VPWR _17246_/B sky130_fd_sc_hd__inv_2
X_13347_ _13310_/A _13347_/B VGND VGND VPWR VPWR _13349_/B sky130_fd_sc_hd__or2_4
X_16135_ _22631_/A VGND VGND VPWR VPWR _16135_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22490__B1 _16918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13278_ _13316_/A _19668_/A VGND VGND VPWR VPWR _13280_/B sky130_fd_sc_hd__or2_4
X_16066_ _24707_/Q VGND VGND VPWR VPWR _16066_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16966__A1_N _24713_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12229_ _25425_/Q VGND VGND VPWR VPWR _12278_/B sky130_fd_sc_hd__inv_2
X_15017_ _24463_/Q VGND VGND VPWR VPWR _15017_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22793__A1 _13593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19825_ _22353_/B _19824_/X _19777_/X _19824_/X VGND VGND VPWR VPWR _23596_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24544__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23284__C _22132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19756_ _19754_/Y _19752_/X _19755_/X _19752_/X VGND VGND VPWR VPWR _23619_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16968_ _24387_/Q VGND VGND VPWR VPWR _17025_/B sky130_fd_sc_hd__inv_2
XANTENNA__21348__A2 _13789_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18707_ _18733_/A VGND VGND VPWR VPWR _18707_/X sky130_fd_sc_hd__buf_2
X_15919_ _15682_/X _15698_/X _15913_/X _15918_/X VGND VGND VPWR VPWR _15920_/A sky130_fd_sc_hd__a211o_4
X_19687_ _13237_/B VGND VGND VPWR VPWR _19687_/Y sky130_fd_sc_hd__inv_2
X_16899_ _22556_/A _16898_/X _16100_/Y _17740_/A VGND VGND VPWR VPWR _16904_/B sky130_fd_sc_hd__a2bb2o_4
X_18638_ _24519_/Q _18757_/A _16611_/Y _18809_/A VGND VGND VPWR VPWR _18638_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18569_ _18566_/A _18572_/B VGND VGND VPWR VPWR _18570_/C sky130_fd_sc_hd__nand2_4
XANTENNA__15983__B1 _15627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16195__A _23232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20600_ _20453_/A _20457_/D _14089_/X VGND VGND VPWR VPWR _23951_/D sky130_fd_sc_hd__o21a_4
XFILLER_36_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21580_ _21580_/A VGND VGND VPWR VPWR _21741_/A sky130_fd_sc_hd__buf_2
XFILLER_21_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20323__A3 _11838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25332__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20531_ _20531_/A _14089_/X _14015_/X VGND VGND VPWR VPWR _20531_/X sky130_fd_sc_hd__and3_4
XANTENNA__22644__B _22644_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23250_ _12864_/A _21872_/X _16916_/Y _22821_/X VGND VGND VPWR VPWR _23250_/X sky130_fd_sc_hd__o22a_4
X_20462_ _14386_/Y _14495_/X _20427_/C VGND VGND VPWR VPWR _20601_/A sky130_fd_sc_hd__a21o_4
X_22201_ _22193_/X _20172_/Y VGND VGND VPWR VPWR _22201_/X sky130_fd_sc_hd__or2_4
XANTENNA__22481__B1 _24712_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23181_ _23181_/A _23101_/B VGND VGND VPWR VPWR _23181_/X sky130_fd_sc_hd__or2_4
X_20393_ _20383_/X _19536_/Y _11867_/A _21200_/A _20380_/X VGND VGND VPWR VPWR _20393_/X
+ sky130_fd_sc_hd__a32o_4
X_22132_ _22132_/A _22132_/B VGND VGND VPWR VPWR _22149_/C sky130_fd_sc_hd__and2_4
XANTENNA__16160__B1 _15474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23025__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22660__A _22660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22063_ _21240_/X VGND VGND VPWR VPWR _22068_/A sky130_fd_sc_hd__buf_2
XFILLER_114_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21014_ _21014_/A _21559_/A _13813_/A _21027_/A VGND VGND VPWR VPWR _21015_/A sky130_fd_sc_hd__or4_4
XFILLER_138_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21276__A _15551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24285__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22536__A1 _17350_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22965_ _22759_/X _22964_/X _22854_/X _12308_/A _22761_/X VGND VGND VPWR VPWR _22966_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_56_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24704_ _24318_/CLK _24704_/D HRESETn VGND VGND VPWR VPWR _24704_/Q sky130_fd_sc_hd__dfrtp_4
X_21916_ _21912_/X _21916_/B _21915_/X VGND VGND VPWR VPWR _21916_/X sky130_fd_sc_hd__and3_4
X_22896_ _22470_/X _22895_/X _21416_/X _12533_/A _22766_/X VGND VGND VPWR VPWR _22897_/B
+ sky130_fd_sc_hd__a32o_4
X_21847_ _12000_/Y _13496_/B _12036_/Y _12072_/D VGND VGND VPWR VPWR _21847_/X sky130_fd_sc_hd__o22a_4
X_24635_ _24654_/CLK _24635_/D HRESETn VGND VGND VPWR VPWR _21322_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15974__B1 _24746_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19165__B1 _19117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _12620_/B _24864_/Q _25398_/Q _12523_/Y VGND VGND VPWR VPWR _12580_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24566_ _24502_/CLK _24566_/D HRESETn VGND VGND VPWR VPWR _16447_/A sky130_fd_sc_hd__dfrtp_4
X_21778_ _19597_/A _21362_/X _23688_/Q _22390_/B VGND VGND VPWR VPWR _21778_/X sky130_fd_sc_hd__o22a_4
XFILLER_93_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22835__A _22835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18425__A1_N _22809_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25073__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20729_ _20728_/Y _20722_/Y _13132_/B VGND VGND VPWR VPWR _20729_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15726__B1 _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23517_ _24309_/CLK _20041_/X VGND VGND VPWR VPWR _20040_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24497_ _24909_/CLK _16641_/X HRESETn VGND VGND VPWR VPWR _23317_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_106_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25002__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _13952_/X _13944_/Y _13959_/Y VGND VGND VPWR VPWR _14251_/D sky130_fd_sc_hd__or3_4
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23448_ _23660_/CLK _23448_/D VGND VGND VPWR VPWR _20221_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23264__A2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ _17453_/A VGND VGND VPWR VPWR _13454_/A sky130_fd_sc_hd__buf_2
XANTENNA__15741__A3 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14181_ _25197_/Q _14181_/B VGND VGND VPWR VPWR _14181_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15449__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23379_ _25098_/CLK _23379_/D VGND VGND VPWR VPWR _23379_/Q sky130_fd_sc_hd__dfxtp_4
X_13132_ _13132_/A _13132_/B VGND VGND VPWR VPWR _13133_/B sky130_fd_sc_hd__or2_4
XFILLER_109_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25118_ _25101_/CLK _25118_/D HRESETn VGND VGND VPWR VPWR _25118_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22570__A _22530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13063_ _13057_/A _13067_/B VGND VGND VPWR VPWR _13063_/Y sky130_fd_sc_hd__nand2_4
X_17940_ _14641_/B _19173_/A VGND VGND VPWR VPWR _17940_/X sky130_fd_sc_hd__or2_4
X_25049_ _23494_/CLK _14754_/X HRESETn VGND VGND VPWR VPWR _14691_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23339__A2_N _24198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18979__B1 _18977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12014_ _12014_/A VGND VGND VPWR VPWR _12014_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17871_ _17874_/A _17867_/X _17871_/C VGND VGND VPWR VPWR _24251_/D sky130_fd_sc_hd__and3_4
Xclkbuf_4_6_0_HCLK clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__13119__D _13119_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19610_ _19609_/X VGND VGND VPWR VPWR _19628_/A sky130_fd_sc_hd__inv_2
X_16822_ _14941_/Y _16819_/X HWDATA[17] _16819_/X VGND VGND VPWR VPWR _16822_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12601__A _12600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19541_ _23691_/Q VGND VGND VPWR VPWR _19541_/Y sky130_fd_sc_hd__inv_2
X_16753_ _16739_/A VGND VGND VPWR VPWR _16753_/X sky130_fd_sc_hd__buf_2
X_13965_ _13917_/X _13965_/B _13964_/X VGND VGND VPWR VPWR _13966_/B sky130_fd_sc_hd__or3_4
XFILLER_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15704_ _15742_/A VGND VGND VPWR VPWR _15713_/A sky130_fd_sc_hd__buf_2
X_12916_ _12850_/B _12915_/X VGND VGND VPWR VPWR _12917_/B sky130_fd_sc_hd__or2_4
X_19472_ _22339_/B _19471_/X _11930_/X _19471_/X VGND VGND VPWR VPWR _23716_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16684_ _16682_/Y _16683_/X _15743_/X _16683_/X VGND VGND VPWR VPWR _16684_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14217__B1 _13800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23937__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13896_ _13895_/X VGND VGND VPWR VPWR _13918_/A sky130_fd_sc_hd__inv_2
XFILLER_62_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18423_ _18396_/X _18404_/X _18413_/X _18422_/X VGND VGND VPWR VPWR _18451_/A sky130_fd_sc_hd__or4_4
X_15635_ _21584_/A _15632_/X _15477_/X _15632_/X VGND VGND VPWR VPWR _24882_/D sky130_fd_sc_hd__a2bb2o_4
X_12847_ _12774_/Y _12833_/Y _12842_/X _12846_/X VGND VGND VPWR VPWR _12847_/X sky130_fd_sc_hd__or4_4
XANTENNA__15965__B1 _15964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19156__B1 _19155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18354_ _17478_/X _17481_/X VGND VGND VPWR VPWR _18355_/A sky130_fd_sc_hd__or2_4
XFILLER_15_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15566_ _15565_/Y _15563_/X _11749_/X _15563_/X VGND VGND VPWR VPWR _24909_/D sky130_fd_sc_hd__a2bb2o_4
X_12778_ _12778_/A VGND VGND VPWR VPWR _12850_/C sky130_fd_sc_hd__inv_2
XFILLER_124_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13789__D _13789_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17305_/A VGND VGND VPWR VPWR _17305_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14517_ _14517_/A VGND VGND VPWR VPWR _14517_/X sky130_fd_sc_hd__buf_2
X_11729_ _15503_/A _15506_/A _11729_/C _11729_/D VGND VGND VPWR VPWR _11730_/D sky130_fd_sc_hd__or4_4
X_18285_ _19492_/B _17725_/X _18278_/D _18319_/B VGND VGND VPWR VPWR _18285_/X sky130_fd_sc_hd__o22a_4
X_15497_ _11719_/B _15494_/X HADDR[20] _15494_/X VGND VGND VPWR VPWR _15497_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12048__A _16183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20710__B1 _20706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17236_ _17236_/A VGND VGND VPWR VPWR _17236_/Y sky130_fd_sc_hd__inv_2
X_14448_ _14436_/Y VGND VGND VPWR VPWR _14448_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16390__B1 _16297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17167_ _16278_/Y _24359_/Q _16278_/Y _24359_/Q VGND VGND VPWR VPWR _17172_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22463__B1 _22447_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24796__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14379_ _14195_/B _18895_/A VGND VGND VPWR VPWR _14394_/B sky130_fd_sc_hd__or2_4
XFILLER_7_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16118_ _16094_/A VGND VGND VPWR VPWR _16118_/X sky130_fd_sc_hd__buf_2
XANTENNA__24725__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17098_ _17007_/Y _17092_/X _17067_/X _17095_/B VGND VGND VPWR VPWR _17099_/A sky130_fd_sc_hd__a211o_4
XANTENNA__22480__A _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_151_0_HCLK clkbuf_7_75_0_HCLK/X VGND VGND VPWR VPWR _24673_/CLK sky130_fd_sc_hd__clkbuf_1
X_16049_ _24713_/Q VGND VGND VPWR VPWR _16049_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19808_ _19802_/Y VGND VGND VPWR VPWR _19808_/X sky130_fd_sc_hd__buf_2
XFILLER_96_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19739_ _13360_/B VGND VGND VPWR VPWR _19739_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19395__B1 _19349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16918__A _16918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22750_ _21580_/A _22750_/B VGND VGND VPWR VPWR _22750_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__14208__B1 _13797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21701_ _24602_/Q _21530_/X VGND VGND VPWR VPWR _21701_/X sky130_fd_sc_hd__or2_4
XFILLER_64_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25513__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15956__B1 _15955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22681_ _22658_/X _22663_/Y _22680_/X VGND VGND VPWR VPWR HRDATA[13] sky130_fd_sc_hd__a21o_4
XANTENNA__21742__A2_N _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19147__B1 _19056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24420_ _24427_/CLK _16820_/X HRESETn VGND VGND VPWR VPWR _14927_/A sky130_fd_sc_hd__dfrtp_4
X_21632_ _21628_/X _21631_/X _14749_/X VGND VGND VPWR VPWR _21632_/X sky130_fd_sc_hd__o21a_4
XANTENNA__13431__B2 _11964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15971__A3 _11803_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24351_ _24355_/CLK _24351_/D HRESETn VGND VGND VPWR VPWR _17237_/A sky130_fd_sc_hd__dfrtp_4
X_21563_ _13511_/Y _21561_/X _12040_/Y _21562_/X VGND VGND VPWR VPWR _21563_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23302_ _21529_/X _23301_/X _23141_/X _24838_/Q _22833_/X VGND VGND VPWR VPWR _23303_/B
+ sky130_fd_sc_hd__a32o_4
X_20514_ _24070_/Q _24075_/Q _20505_/C VGND VGND VPWR VPWR _20515_/D sky130_fd_sc_hd__or3_4
X_24282_ _24278_/CLK _24282_/D HRESETn VGND VGND VPWR VPWR _17576_/A sky130_fd_sc_hd__dfrtp_4
X_21494_ _21469_/X _21491_/X _21493_/X VGND VGND VPWR VPWR _21494_/Y sky130_fd_sc_hd__a21oi_4
X_23233_ _16469_/A _23166_/X _23130_/X VGND VGND VPWR VPWR _23233_/X sky130_fd_sc_hd__o21a_4
X_20445_ _20496_/C _20445_/B _20422_/Y VGND VGND VPWR VPWR _20446_/B sky130_fd_sc_hd__and3_4
XFILLER_107_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24466__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23164_ _23128_/A _23163_/X VGND VGND VPWR VPWR _23176_/B sky130_fd_sc_hd__nor2_4
X_20376_ _20375_/Y _20373_/X _19632_/A _20373_/X VGND VGND VPWR VPWR _23389_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12405__B _13008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22115_ _22114_/X VGND VGND VPWR VPWR _22115_/Y sky130_fd_sc_hd__inv_2
X_23095_ _21108_/B VGND VGND VPWR VPWR _23095_/X sky130_fd_sc_hd__buf_2
XFILLER_88_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14695__B1 _21612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22046_ _22046_/A _19585_/A VGND VGND VPWR VPWR _22046_/X sky130_fd_sc_hd__and2_4
XFILLER_125_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21734__A _16533_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23997_ _24885_/CLK _23997_/D HRESETn VGND VGND VPWR VPWR _23997_/Q sky130_fd_sc_hd__dfrtp_4
X_13750_ _13757_/B VGND VGND VPWR VPWR _13751_/A sky130_fd_sc_hd__inv_2
XFILLER_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22948_ _22948_/A VGND VGND VPWR VPWR _22948_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25254__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12701_ _12529_/Y _12665_/A VGND VGND VPWR VPWR _12735_/A sky130_fd_sc_hd__or2_4
XFILLER_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13681_ _11682_/Y _11689_/Y VGND VGND VPWR VPWR _13729_/B sky130_fd_sc_hd__or2_4
XANTENNA__15947__B1 _24761_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19138__B1 _19136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_14_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22879_ _22879_/A VGND VGND VPWR VPWR _22879_/X sky130_fd_sc_hd__buf_2
X_15420_ _15415_/X _15419_/Y _15407_/X VGND VGND VPWR VPWR _24965_/D sky130_fd_sc_hd__and3_4
XFILLER_19_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13252__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12632_ _12632_/A VGND VGND VPWR VPWR _12632_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24618_ _24346_/CLK _24618_/D HRESETn VGND VGND VPWR VPWR _22899_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12225__A2 _21526_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22565__A _21009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _24847_/Q VGND VGND VPWR VPWR _12563_/Y sky130_fd_sc_hd__inv_2
X_15351_ _15336_/A _15336_/B VGND VGND VPWR VPWR _15352_/B sky130_fd_sc_hd__or2_4
XFILLER_15_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24549_ _24465_/CLK _16502_/X HRESETn VGND VGND VPWR VPWR _16501_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22284__B _21073_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14302_ _14299_/Y VGND VGND VPWR VPWR _14302_/X sky130_fd_sc_hd__buf_2
X_18070_ _17982_/X _23737_/Q VGND VGND VPWR VPWR _18070_/X sky130_fd_sc_hd__or2_4
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _25425_/Q _12494_/B VGND VGND VPWR VPWR _12494_/X sky130_fd_sc_hd__or2_4
X_15282_ _15282_/A _15282_/B _15281_/Y VGND VGND VPWR VPWR _24997_/D sky130_fd_sc_hd__and3_4
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23237__A2 _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17021_ _17020_/X VGND VGND VPWR VPWR _17064_/A sky130_fd_sc_hd__buf_2
X_14233_ _25184_/Q VGND VGND VPWR VPWR _14233_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22445__B1 _16603_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14164_ _14125_/A _14163_/Y _14099_/A _14125_/A VGND VGND VPWR VPWR _25201_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13115_ _13106_/X _13115_/B _13115_/C VGND VGND VPWR VPWR _25323_/D sky130_fd_sc_hd__and3_4
XFILLER_3_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24136__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_224_0_HCLK clkbuf_8_225_0_HCLK/A VGND VGND VPWR VPWR _25374_/CLK sky130_fd_sc_hd__clkbuf_1
X_14095_ _20977_/B VGND VGND VPWR VPWR _20978_/B sky130_fd_sc_hd__inv_2
X_18972_ _18972_/A VGND VGND VPWR VPWR _18972_/X sky130_fd_sc_hd__buf_2
XFILLER_98_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13046_ _13048_/B VGND VGND VPWR VPWR _13047_/B sky130_fd_sc_hd__inv_2
X_17923_ _17920_/B _17920_/C VGND VGND VPWR VPWR _17923_/X sky130_fd_sc_hd__or2_4
XFILLER_79_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21420__A1 _21413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17854_ _17744_/Y _17854_/B VGND VGND VPWR VPWR _17855_/C sky130_fd_sc_hd__or2_4
XFILLER_113_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12331__A _24816_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16805_ _14905_/Y _16802_/X HWDATA[27] _16802_/X VGND VGND VPWR VPWR _16805_/X sky130_fd_sc_hd__a2bb2o_4
X_17785_ _17785_/A _17790_/B VGND VGND VPWR VPWR _17787_/B sky130_fd_sc_hd__or2_4
XFILLER_54_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14989__B2 _24448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14997_ _15197_/A _24458_/Q _15197_/A _24458_/Q VGND VGND VPWR VPWR _15002_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19524_ _19523_/Y _19521_/X _11943_/X _19521_/X VGND VGND VPWR VPWR _19524_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15642__A _15642_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16736_ _24461_/Q VGND VGND VPWR VPWR _16736_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13948_ _13935_/D VGND VGND VPWR VPWR _13948_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_1_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19455_ _19454_/Y _19452_/X _19364_/X _19452_/X VGND VGND VPWR VPWR _23721_/D sky130_fd_sc_hd__a2bb2o_4
X_16667_ _16666_/Y _16664_/X _16398_/X _16664_/X VGND VGND VPWR VPWR _24488_/D sky130_fd_sc_hd__a2bb2o_4
X_13879_ _13871_/X _13878_/X _25174_/Q _13856_/Y VGND VGND VPWR VPWR _13879_/X sky130_fd_sc_hd__o22a_4
X_18406_ _16216_/A _24164_/Q _16216_/Y _18405_/Y VGND VGND VPWR VPWR _18413_/A sky130_fd_sc_hd__o22a_4
XFILLER_90_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13162__A _13162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15618_ _15616_/Y _15612_/X _11829_/X _15617_/X VGND VGND VPWR VPWR _24888_/D sky130_fd_sc_hd__a2bb2o_4
X_19386_ _23745_/Q VGND VGND VPWR VPWR _19386_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16598_ _16597_/Y _16595_/X _16340_/X _16595_/X VGND VGND VPWR VPWR _16598_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22475__A _22419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18337_ _17459_/X _17451_/Y _18335_/X VGND VGND VPWR VPWR _18337_/X sky130_fd_sc_hd__o21a_4
X_15549_ _15549_/A _15549_/B VGND VGND VPWR VPWR _15549_/X sky130_fd_sc_hd__or2_4
XANTENNA__17569__A _17630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24977__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16473__A _24560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18268_ _13795_/D _18253_/X _18267_/X _24209_/Q _18262_/A VGND VGND VPWR VPWR _18268_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24906__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17219_ _16354_/Y _24332_/Q _24627_/Q _17234_/A VGND VGND VPWR VPWR _17224_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22487__A2_N _22482_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22436__B1 _25363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19784__A _19793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18199_ _17982_/X _23765_/Q VGND VGND VPWR VPWR _18199_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_34_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_69_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12506__A _13008_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20230_ _13183_/B VGND VGND VPWR VPWR _20230_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19522__A2_N _19516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20161_ _20161_/A VGND VGND VPWR VPWR _20161_/X sky130_fd_sc_hd__buf_2
XFILLER_103_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15817__A _15817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14721__A _14705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17735__C _24198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20092_ _20092_/A VGND VGND VPWR VPWR _20092_/X sky130_fd_sc_hd__buf_2
XFILLER_135_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23920_ _24945_/CLK _23920_/D HRESETn VGND VGND VPWR VPWR _23920_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14429__B1 _14239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23851_ _24398_/CLK _19089_/X VGND VGND VPWR VPWR _23851_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22802_ _16223_/A _22884_/B VGND VGND VPWR VPWR _22802_/X sky130_fd_sc_hd__or2_4
X_20994_ _23968_/D VGND VGND VPWR VPWR _20996_/A sky130_fd_sc_hd__inv_2
XFILLER_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23782_ _23846_/CLK _19281_/X VGND VGND VPWR VPWR _23782_/Q sky130_fd_sc_hd__dfxtp_4
X_25521_ _24275_/CLK _11806_/X HRESETn VGND VGND VPWR VPWR _11802_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22733_ _22733_/A _22522_/B VGND VGND VPWR VPWR _22736_/B sky130_fd_sc_hd__or2_4
XFILLER_111_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25452_ _24383_/CLK _12176_/X HRESETn VGND VGND VPWR VPWR _25452_/Q sky130_fd_sc_hd__dfrtp_4
X_22664_ _15019_/Y _22664_/B VGND VGND VPWR VPWR _22664_/X sky130_fd_sc_hd__and2_4
XFILLER_40_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21615_ _14680_/X VGND VGND VPWR VPWR _21616_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_116_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_233_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24403_ _24435_/CLK _16853_/X HRESETn VGND VGND VPWR VPWR _24403_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22816__C _22493_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25383_ _25385_/CLK _12876_/Y HRESETn VGND VGND VPWR VPWR _25383_/Q sky130_fd_sc_hd__dfrtp_4
X_22595_ _22595_/A _21085_/A VGND VGND VPWR VPWR _22595_/X sky130_fd_sc_hd__or2_4
XFILLER_55_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19540__B1 _19426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13800__A _16359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21546_ _21331_/X _21545_/X VGND VGND VPWR VPWR _21546_/Y sky130_fd_sc_hd__nor2_4
XFILLER_90_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24647__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24334_ _24334_/CLK _17370_/X HRESETn VGND VGND VPWR VPWR _17168_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_127_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22427__B1 _11828_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24265_ _24692_/CLK _17817_/Y HRESETn VGND VGND VPWR VPWR _16941_/A sky130_fd_sc_hd__dfrtp_4
X_21477_ _21477_/A _19904_/Y VGND VGND VPWR VPWR _21480_/B sky130_fd_sc_hd__or2_4
XANTENNA__12416__A _12277_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22832__B _22832_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23216_ _24627_/Q _21519_/B VGND VGND VPWR VPWR _23216_/X sky130_fd_sc_hd__or2_4
X_20428_ _13976_/X _20428_/B _20428_/C _20428_/D VGND VGND VPWR VPWR _20428_/X sky130_fd_sc_hd__or4_4
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21729__A _21729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24196_ _24187_/CLK _18332_/X HRESETn VGND VGND VPWR VPWR _24196_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23147_ _16295_/A _22898_/X VGND VGND VPWR VPWR _23147_/X sky130_fd_sc_hd__or2_4
X_20359_ _18275_/A _19971_/X _19492_/X VGND VGND VPWR VPWR _20360_/A sky130_fd_sc_hd__or3_4
XFILLER_49_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23366__D scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23078_ _24053_/Q _21287_/Y _24021_/Q _21589_/X VGND VGND VPWR VPWR _23078_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_66_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14920_ _25019_/Q _14919_/A _15194_/A _14919_/Y VGND VGND VPWR VPWR _14920_/X sky130_fd_sc_hd__o22a_4
X_22029_ _22024_/A _22029_/B VGND VGND VPWR VPWR _22029_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_54_0_HCLK clkbuf_8_55_0_HCLK/A VGND VGND VPWR VPWR _24376_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_48_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25435__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14851_ _14843_/X _14850_/Y _14815_/C _14843_/X VGND VGND VPWR VPWR _14851_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22279__B _22406_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19359__B1 _19291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13802_ _13802_/A VGND VGND VPWR VPWR _13802_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17570_ _24291_/Q VGND VGND VPWR VPWR _17580_/A sky130_fd_sc_hd__inv_2
X_14782_ _14781_/X VGND VGND VPWR VPWR _16880_/A sky130_fd_sc_hd__buf_2
X_11994_ _11994_/A _11994_/B VGND VGND VPWR VPWR _11994_/X sky130_fd_sc_hd__and2_4
XFILLER_21_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14840__B1 _25184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16521_ _16057_/A VGND VGND VPWR VPWR _16521_/X sky130_fd_sc_hd__buf_2
X_13733_ _25268_/Q _13721_/X _13703_/X _11689_/Y VGND VGND VPWR VPWR _13733_/X sky130_fd_sc_hd__o22a_4
XFILLER_56_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19240_ _19239_/Y _19235_/X _19149_/X _19221_/Y VGND VGND VPWR VPWR _19240_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16452_ _16452_/A VGND VGND VPWR VPWR _22736_/A sky130_fd_sc_hd__buf_2
XFILLER_31_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15396__A1 _15073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14199__A2 _14196_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13664_ _13664_/A _13650_/X _20900_/A VGND VGND VPWR VPWR _13664_/X sky130_fd_sc_hd__or3_4
XANTENNA__16593__B1 _16238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15403_ _15384_/A _15400_/B _15403_/C VGND VGND VPWR VPWR _24971_/D sky130_fd_sc_hd__and3_4
X_12615_ _25389_/Q VGND VGND VPWR VPWR _12728_/A sky130_fd_sc_hd__inv_2
X_19171_ _18219_/B VGND VGND VPWR VPWR _19171_/Y sky130_fd_sc_hd__inv_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16383_ _15109_/Y _16375_/X _16380_/X _16382_/X VGND VGND VPWR VPWR _24596_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ _13595_/A VGND VGND VPWR VPWR _13815_/A sky130_fd_sc_hd__buf_2
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18122_ _18186_/A _18122_/B VGND VGND VPWR VPWR _18124_/B sky130_fd_sc_hd__or2_4
XANTENNA__19531__B1 _11955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15334_ _15315_/A _15329_/Y _15333_/X VGND VGND VPWR VPWR _15334_/X sky130_fd_sc_hd__or3_4
XANTENNA__24388__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12546_ _24871_/Q VGND VGND VPWR VPWR _12546_/Y sky130_fd_sc_hd__inv_2
X_18053_ _18184_/A _18053_/B _18053_/C VGND VGND VPWR VPWR _18058_/B sky130_fd_sc_hd__and3_4
XANTENNA__24317__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15265_ _15265_/A VGND VGND VPWR VPWR _25003_/D sky130_fd_sc_hd__inv_2
X_12477_ _12220_/X _12203_/X _12471_/X VGND VGND VPWR VPWR _12477_/X sky130_fd_sc_hd__or3_4
X_17004_ _16019_/Y _24382_/Q _24713_/Q _17041_/D VGND VGND VPWR VPWR _17004_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22742__B _22592_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14216_ _20664_/A VGND VGND VPWR VPWR _14216_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15196_ _25020_/Q _15195_/Y VGND VGND VPWR VPWR _15196_/X sky130_fd_sc_hd__or2_4
XFILLER_98_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14147_ _14116_/A _14116_/B _14116_/A _14116_/B VGND VGND VPWR VPWR _14147_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_28_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14078_ _14078_/A VGND VGND VPWR VPWR _14078_/X sky130_fd_sc_hd__buf_2
X_18955_ _16781_/X VGND VGND VPWR VPWR _18955_/X sky130_fd_sc_hd__buf_2
XANTENNA__13157__A _13156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13029_ _13029_/A _13029_/B VGND VGND VPWR VPWR _13038_/B sky130_fd_sc_hd__or2_4
X_17906_ _17898_/Y _17905_/A _17904_/X _24243_/Q _17905_/Y VGND VGND VPWR VPWR _24243_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18886_ _20582_/B VGND VGND VPWR VPWR _18886_/X sky130_fd_sc_hd__buf_2
XANTENNA__23952__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17837_ _17837_/A _17751_/X VGND VGND VPWR VPWR _17837_/X sky130_fd_sc_hd__or2_4
XANTENNA__25105__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17768_ _23314_/A _17768_/B VGND VGND VPWR VPWR _17768_/Y sky130_fd_sc_hd__nand2_4
XFILLER_82_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16719_ _16719_/A VGND VGND VPWR VPWR _16719_/Y sky130_fd_sc_hd__inv_2
X_19507_ _19494_/Y VGND VGND VPWR VPWR _19507_/X sky130_fd_sc_hd__buf_2
XANTENNA__13604__B _13610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17699_ _17699_/A VGND VGND VPWR VPWR _17699_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19438_ _19431_/A VGND VGND VPWR VPWR _19438_/X sky130_fd_sc_hd__buf_2
XFILLER_74_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16584__B1 _16325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19369_ _19355_/Y VGND VGND VPWR VPWR _19369_/X sky130_fd_sc_hd__buf_2
XANTENNA__22657__B1 _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21400_ _21385_/A _20098_/Y VGND VGND VPWR VPWR _21400_/X sky130_fd_sc_hd__or2_4
XFILLER_124_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22380_ _14716_/A _22359_/Y _22366_/Y _22373_/Y _22379_/Y VGND VGND VPWR VPWR _22380_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24740__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21331_ _21331_/A VGND VGND VPWR VPWR _21331_/X sky130_fd_sc_hd__buf_2
XANTENNA__24058__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15160__A2_N _15077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24050_ _24487_/CLK _24050_/D HRESETn VGND VGND VPWR VPWR _24050_/Q sky130_fd_sc_hd__dfrtp_4
X_21262_ _13817_/A VGND VGND VPWR VPWR _22575_/A sky130_fd_sc_hd__buf_2
XFILLER_128_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19825__B2 _19824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23001_ _23065_/A _23001_/B _23000_/X VGND VGND VPWR VPWR _23002_/D sky130_fd_sc_hd__and3_4
X_20213_ _20209_/Y _20212_/X _18247_/X _20212_/X VGND VGND VPWR VPWR _23452_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15547__A _22873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21193_ _21185_/A _19947_/Y VGND VGND VPWR VPWR _21194_/C sky130_fd_sc_hd__or2_4
XFILLER_85_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20144_ _20144_/A VGND VGND VPWR VPWR _20144_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19589__B1 _19426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20075_ _20065_/A _18325_/X _11867_/A _23501_/Q _20065_/Y VGND VGND VPWR VPWR _20075_/X
+ sky130_fd_sc_hd__a32o_4
X_24952_ _24950_/CLK _15453_/X HRESETn VGND VGND VPWR VPWR _24952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23903_ _24209_/CLK _23903_/D VGND VGND VPWR VPWR _13379_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17481__B _17449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24883_ _24883_/CLK _15633_/X HRESETn VGND VGND VPWR VPWR _24883_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23834_ _23826_/CLK _23834_/D VGND VGND VPWR VPWR _23834_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_113_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21148__B1 _14190_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20977_ _20978_/A _20977_/B _20977_/C VGND VGND VPWR VPWR _20977_/X sky130_fd_sc_hd__and3_4
XANTENNA__22896__B1 _12533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24899__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23765_ _23772_/CLK _23765_/D VGND VGND VPWR VPWR _23765_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25504_ _25503_/CLK _11898_/X HRESETn VGND VGND VPWR VPWR _11869_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__24828__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22716_ _22716_/A VGND VGND VPWR VPWR _22716_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23696_ _24930_/CLK _19526_/X VGND VGND VPWR VPWR _23696_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23004__A _23004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22648__B1 _24820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25435_ _25449_/CLK _25435_/D HRESETn VGND VGND VPWR VPWR _12248_/A sky130_fd_sc_hd__dfrtp_4
X_22647_ _24748_/Q _22644_/B VGND VGND VPWR VPWR _22647_/X sky130_fd_sc_hd__or2_4
XANTENNA__18316__A1 _18298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22112__A2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12400_ _12385_/A _12398_/A VGND VGND VPWR VPWR _12400_/X sky130_fd_sc_hd__or2_4
X_13380_ _13312_/A _23503_/Q VGND VGND VPWR VPWR _13381_/C sky130_fd_sc_hd__or2_4
XFILLER_55_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24481__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25366_ _25330_/CLK _25366_/D HRESETn VGND VGND VPWR VPWR _25366_/Q sky130_fd_sc_hd__dfrtp_4
X_22578_ _22505_/X _22576_/X _21950_/X _22577_/X VGND VGND VPWR VPWR _22578_/X sky130_fd_sc_hd__o22a_4
XFILLER_127_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22843__A _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12331_ _24816_/Q VGND VGND VPWR VPWR _12331_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24410__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24317_ _24883_/CLK _24317_/D HRESETn VGND VGND VPWR VPWR _24317_/Q sky130_fd_sc_hd__dfrtp_4
X_21529_ _21108_/B VGND VGND VPWR VPWR _21529_/X sky130_fd_sc_hd__buf_2
X_25297_ _25301_/CLK _13510_/X HRESETn VGND VGND VPWR VPWR _13509_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14889__B1 _14888_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12262_ _12253_/X _12262_/B _12258_/X _12261_/X VGND VGND VPWR VPWR _12262_/X sky130_fd_sc_hd__or4_4
X_15050_ _15071_/A _24459_/Q _15212_/A _24453_/Q VGND VGND VPWR VPWR _15054_/C sky130_fd_sc_hd__a2bb2o_4
X_24248_ _24248_/CLK _17880_/X HRESETn VGND VGND VPWR VPWR _24248_/Q sky130_fd_sc_hd__dfrtp_4
X_14001_ _14001_/A _13989_/A _13999_/X _14001_/D VGND VGND VPWR VPWR _14001_/X sky130_fd_sc_hd__or4_4
XFILLER_108_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12193_ _22964_/A VGND VGND VPWR VPWR _12193_/Y sky130_fd_sc_hd__inv_2
X_24179_ _23933_/CLK _18387_/X HRESETn VGND VGND VPWR VPWR _24179_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18740_ _18733_/A _18737_/B _18740_/C VGND VGND VPWR VPWR _18740_/X sky130_fd_sc_hd__or3_4
XFILLER_114_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15952_ HWDATA[22] VGND VGND VPWR VPWR _15952_/X sky130_fd_sc_hd__buf_2
XFILLER_103_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14903_ _15065_/A VGND VGND VPWR VPWR _14903_/X sky130_fd_sc_hd__buf_2
XFILLER_49_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18671_ _18671_/A VGND VGND VPWR VPWR _18698_/C sky130_fd_sc_hd__inv_2
X_15883_ _12779_/Y _15879_/X _11784_/X _15882_/X VGND VGND VPWR VPWR _15883_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17622_ _17885_/B _17618_/Y _17621_/X VGND VGND VPWR VPWR _17623_/A sky130_fd_sc_hd__or3_4
X_14834_ _14817_/C _14803_/B _14817_/C _14803_/B VGND VGND VPWR VPWR _14834_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13077__C1 _13031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17553_ _17792_/C VGND VGND VPWR VPWR _17837_/A sky130_fd_sc_hd__buf_2
X_14765_ _13738_/A VGND VGND VPWR VPWR _16173_/A sky130_fd_sc_hd__buf_2
XANTENNA__19599__A _18254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22887__B1 _22524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11977_ _11972_/X _11976_/X VGND VGND VPWR VPWR _11977_/X sky130_fd_sc_hd__and2_4
X_16504_ _16504_/A VGND VGND VPWR VPWR _16504_/X sky130_fd_sc_hd__buf_2
XFILLER_45_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13716_ _11685_/Y _13688_/B VGND VGND VPWR VPWR _13716_/Y sky130_fd_sc_hd__nand2_4
X_17484_ _17483_/X VGND VGND VPWR VPWR _17484_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16566__B1 _16306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24569__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14696_ _14719_/B VGND VGND VPWR VPWR _14698_/C sky130_fd_sc_hd__inv_2
XFILLER_108_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19223_ _19218_/Y _19222_/X _19155_/X _19222_/X VGND VGND VPWR VPWR _19223_/X sky130_fd_sc_hd__a2bb2o_4
X_16435_ _15126_/Y _16433_/X _16064_/X _16433_/X VGND VGND VPWR VPWR _16435_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22639__B1 _12235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13647_ _25287_/Q _13640_/X _24084_/D VGND VGND VPWR VPWR _25287_/D sky130_fd_sc_hd__o21a_4
XFILLER_73_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19154_ _19153_/Y VGND VGND VPWR VPWR _19154_/X sky130_fd_sc_hd__buf_2
XFILLER_73_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16366_ _16720_/A VGND VGND VPWR VPWR _16366_/X sky130_fd_sc_hd__buf_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _13567_/X _13578_/B _13574_/X _13578_/D VGND VGND VPWR VPWR _13578_/X sky130_fd_sc_hd__or4_4
XFILLER_34_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18105_ _18137_/A _18103_/X _18105_/C VGND VGND VPWR VPWR _18106_/C sky130_fd_sc_hd__and3_4
X_15317_ _15309_/X _15316_/X _15155_/Y VGND VGND VPWR VPWR _15317_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12529_ _25388_/Q VGND VGND VPWR VPWR _12529_/Y sky130_fd_sc_hd__inv_2
X_19085_ _19084_/X VGND VGND VPWR VPWR _19098_/A sky130_fd_sc_hd__inv_2
X_16297_ HWDATA[26] VGND VGND VPWR VPWR _16297_/X sky130_fd_sc_hd__buf_2
XFILLER_9_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18036_ _18211_/A _18036_/B VGND VGND VPWR VPWR _18036_/X sky130_fd_sc_hd__or2_4
X_15248_ _15248_/A _15248_/B VGND VGND VPWR VPWR _15249_/B sky130_fd_sc_hd__or2_4
XANTENNA__23064__B1 _22997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15541__B2 _15538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12355__B2 _24830_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15179_ _15179_/A _15179_/B VGND VGND VPWR VPWR _15181_/B sky130_fd_sc_hd__or2_4
XFILLER_113_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25357__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19987_ _19987_/A VGND VGND VPWR VPWR _21804_/B sky130_fd_sc_hd__inv_2
XFILLER_80_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18938_ _18936_/Y _18937_/X _16852_/X _18937_/X VGND VGND VPWR VPWR _23903_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21816__B _21816_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

