magic
tech sky130A
magscale 1 2
timestamp 1609333376
<< obsli1 >>
rect 1104 1879 119019 77529
<< obsm1 >>
rect 1104 1848 119034 77640
<< obsm2 >>
rect 1398 23 119122 79385
<< metal3 >>
rect 0 79152 800 79272
rect 119200 79288 120000 79408
rect 119200 78608 120000 78728
rect 0 78200 800 78320
rect 119200 78064 120000 78184
rect 0 77248 800 77368
rect 119200 77384 120000 77504
rect 119200 76840 120000 76960
rect 0 76296 800 76416
rect 119200 76160 120000 76280
rect 0 75344 800 75464
rect 119200 75480 120000 75600
rect 119200 74936 120000 75056
rect 0 74392 800 74512
rect 119200 74256 120000 74376
rect 119200 73712 120000 73832
rect 0 73440 800 73560
rect 119200 73032 120000 73152
rect 0 72488 800 72608
rect 119200 72352 120000 72472
rect 119200 71808 120000 71928
rect 0 71536 800 71656
rect 119200 71128 120000 71248
rect 0 70584 800 70704
rect 119200 70584 120000 70704
rect 119200 69904 120000 70024
rect 0 69632 800 69752
rect 119200 69224 120000 69344
rect 0 68680 800 68800
rect 119200 68680 120000 68800
rect 119200 68000 120000 68120
rect 0 67728 800 67848
rect 119200 67456 120000 67576
rect 0 66776 800 66896
rect 119200 66776 120000 66896
rect 119200 66096 120000 66216
rect 0 65824 800 65944
rect 119200 65552 120000 65672
rect 0 64872 800 64992
rect 119200 64872 120000 64992
rect 119200 64328 120000 64448
rect 0 63920 800 64040
rect 119200 63648 120000 63768
rect 0 62968 800 63088
rect 119200 62968 120000 63088
rect 119200 62424 120000 62544
rect 0 62016 800 62136
rect 119200 61744 120000 61864
rect 0 61064 800 61184
rect 119200 61200 120000 61320
rect 119200 60520 120000 60640
rect 0 60112 800 60232
rect 119200 59976 120000 60096
rect 0 59160 800 59280
rect 119200 59296 120000 59416
rect 119200 58616 120000 58736
rect 0 58208 800 58328
rect 119200 58072 120000 58192
rect 0 57256 800 57376
rect 119200 57392 120000 57512
rect 119200 56848 120000 56968
rect 0 56304 800 56424
rect 119200 56168 120000 56288
rect 0 55352 800 55472
rect 119200 55488 120000 55608
rect 119200 54944 120000 55064
rect 0 54400 800 54520
rect 119200 54264 120000 54384
rect 119200 53720 120000 53840
rect 0 53448 800 53568
rect 119200 53040 120000 53160
rect 0 52496 800 52616
rect 119200 52360 120000 52480
rect 119200 51816 120000 51936
rect 0 51544 800 51664
rect 119200 51136 120000 51256
rect 0 50592 800 50712
rect 119200 50592 120000 50712
rect 119200 49912 120000 50032
rect 0 49640 800 49760
rect 119200 49232 120000 49352
rect 0 48688 800 48808
rect 119200 48688 120000 48808
rect 119200 48008 120000 48128
rect 0 47736 800 47856
rect 119200 47464 120000 47584
rect 0 46784 800 46904
rect 119200 46784 120000 46904
rect 119200 46104 120000 46224
rect 0 45832 800 45952
rect 119200 45560 120000 45680
rect 0 44880 800 45000
rect 119200 44880 120000 45000
rect 119200 44336 120000 44456
rect 0 43928 800 44048
rect 119200 43656 120000 43776
rect 0 42976 800 43096
rect 119200 42976 120000 43096
rect 119200 42432 120000 42552
rect 0 42024 800 42144
rect 119200 41752 120000 41872
rect 0 41072 800 41192
rect 119200 41208 120000 41328
rect 119200 40528 120000 40648
rect 0 40120 800 40240
rect 119200 39984 120000 40104
rect 0 39168 800 39288
rect 119200 39304 120000 39424
rect 119200 38624 120000 38744
rect 0 38216 800 38336
rect 119200 38080 120000 38200
rect 0 37264 800 37384
rect 119200 37400 120000 37520
rect 119200 36856 120000 36976
rect 0 36312 800 36432
rect 119200 36176 120000 36296
rect 0 35360 800 35480
rect 119200 35496 120000 35616
rect 119200 34952 120000 35072
rect 0 34408 800 34528
rect 119200 34272 120000 34392
rect 119200 33728 120000 33848
rect 0 33456 800 33576
rect 119200 33048 120000 33168
rect 0 32504 800 32624
rect 119200 32368 120000 32488
rect 119200 31824 120000 31944
rect 0 31552 800 31672
rect 119200 31144 120000 31264
rect 0 30600 800 30720
rect 119200 30600 120000 30720
rect 119200 29920 120000 30040
rect 0 29648 800 29768
rect 119200 29240 120000 29360
rect 0 28696 800 28816
rect 119200 28696 120000 28816
rect 119200 28016 120000 28136
rect 0 27744 800 27864
rect 119200 27472 120000 27592
rect 0 26792 800 26912
rect 119200 26792 120000 26912
rect 119200 26112 120000 26232
rect 0 25840 800 25960
rect 119200 25568 120000 25688
rect 0 24888 800 25008
rect 119200 24888 120000 25008
rect 119200 24344 120000 24464
rect 0 23936 800 24056
rect 119200 23664 120000 23784
rect 0 22984 800 23104
rect 119200 22984 120000 23104
rect 119200 22440 120000 22560
rect 0 22032 800 22152
rect 119200 21760 120000 21880
rect 0 21080 800 21200
rect 119200 21216 120000 21336
rect 119200 20536 120000 20656
rect 0 20128 800 20248
rect 119200 19992 120000 20112
rect 0 19176 800 19296
rect 119200 19312 120000 19432
rect 119200 18632 120000 18752
rect 0 18224 800 18344
rect 119200 18088 120000 18208
rect 0 17272 800 17392
rect 119200 17408 120000 17528
rect 119200 16864 120000 16984
rect 0 16320 800 16440
rect 119200 16184 120000 16304
rect 0 15368 800 15488
rect 119200 15504 120000 15624
rect 119200 14960 120000 15080
rect 0 14416 800 14536
rect 119200 14280 120000 14400
rect 119200 13736 120000 13856
rect 0 13464 800 13584
rect 119200 13056 120000 13176
rect 0 12512 800 12632
rect 119200 12376 120000 12496
rect 119200 11832 120000 11952
rect 0 11560 800 11680
rect 119200 11152 120000 11272
rect 0 10608 800 10728
rect 119200 10608 120000 10728
rect 119200 9928 120000 10048
rect 0 9656 800 9776
rect 119200 9248 120000 9368
rect 0 8704 800 8824
rect 119200 8704 120000 8824
rect 119200 8024 120000 8144
rect 0 7752 800 7872
rect 119200 7480 120000 7600
rect 0 6800 800 6920
rect 119200 6800 120000 6920
rect 119200 6120 120000 6240
rect 0 5848 800 5968
rect 119200 5576 120000 5696
rect 0 4896 800 5016
rect 119200 4896 120000 5016
rect 119200 4352 120000 4472
rect 0 3944 800 4064
rect 119200 3672 120000 3792
rect 0 2992 800 3112
rect 119200 2992 120000 3112
rect 119200 2448 120000 2568
rect 0 2040 800 2160
rect 119200 1768 120000 1888
rect 0 1088 800 1208
rect 119200 1224 120000 1344
rect 119200 544 120000 664
rect 0 136 800 256
rect 119200 0 120000 120
<< obsm3 >>
rect 800 79352 119120 79381
rect 880 79208 119120 79352
rect 880 79072 119200 79208
rect 800 78808 119200 79072
rect 800 78528 119120 78808
rect 800 78400 119200 78528
rect 880 78264 119200 78400
rect 880 78120 119120 78264
rect 800 77984 119120 78120
rect 800 77584 119200 77984
rect 800 77448 119120 77584
rect 880 77304 119120 77448
rect 880 77168 119200 77304
rect 800 77040 119200 77168
rect 800 76760 119120 77040
rect 800 76496 119200 76760
rect 880 76360 119200 76496
rect 880 76216 119120 76360
rect 800 76080 119120 76216
rect 800 75680 119200 76080
rect 800 75544 119120 75680
rect 880 75400 119120 75544
rect 880 75264 119200 75400
rect 800 75136 119200 75264
rect 800 74856 119120 75136
rect 800 74592 119200 74856
rect 880 74456 119200 74592
rect 880 74312 119120 74456
rect 800 74176 119120 74312
rect 800 73912 119200 74176
rect 800 73640 119120 73912
rect 880 73632 119120 73640
rect 880 73360 119200 73632
rect 800 73232 119200 73360
rect 800 72952 119120 73232
rect 800 72688 119200 72952
rect 880 72552 119200 72688
rect 880 72408 119120 72552
rect 800 72272 119120 72408
rect 800 72008 119200 72272
rect 800 71736 119120 72008
rect 880 71728 119120 71736
rect 880 71456 119200 71728
rect 800 71328 119200 71456
rect 800 71048 119120 71328
rect 800 70784 119200 71048
rect 880 70504 119120 70784
rect 800 70104 119200 70504
rect 800 69832 119120 70104
rect 880 69824 119120 69832
rect 880 69552 119200 69824
rect 800 69424 119200 69552
rect 800 69144 119120 69424
rect 800 68880 119200 69144
rect 880 68600 119120 68880
rect 800 68200 119200 68600
rect 800 67928 119120 68200
rect 880 67920 119120 67928
rect 880 67656 119200 67920
rect 880 67648 119120 67656
rect 800 67376 119120 67648
rect 800 66976 119200 67376
rect 880 66696 119120 66976
rect 800 66296 119200 66696
rect 800 66024 119120 66296
rect 880 66016 119120 66024
rect 880 65752 119200 66016
rect 880 65744 119120 65752
rect 800 65472 119120 65744
rect 800 65072 119200 65472
rect 880 64792 119120 65072
rect 800 64528 119200 64792
rect 800 64248 119120 64528
rect 800 64120 119200 64248
rect 880 63848 119200 64120
rect 880 63840 119120 63848
rect 800 63568 119120 63840
rect 800 63168 119200 63568
rect 880 62888 119120 63168
rect 800 62624 119200 62888
rect 800 62344 119120 62624
rect 800 62216 119200 62344
rect 880 61944 119200 62216
rect 880 61936 119120 61944
rect 800 61664 119120 61936
rect 800 61400 119200 61664
rect 800 61264 119120 61400
rect 880 61120 119120 61264
rect 880 60984 119200 61120
rect 800 60720 119200 60984
rect 800 60440 119120 60720
rect 800 60312 119200 60440
rect 880 60176 119200 60312
rect 880 60032 119120 60176
rect 800 59896 119120 60032
rect 800 59496 119200 59896
rect 800 59360 119120 59496
rect 880 59216 119120 59360
rect 880 59080 119200 59216
rect 800 58816 119200 59080
rect 800 58536 119120 58816
rect 800 58408 119200 58536
rect 880 58272 119200 58408
rect 880 58128 119120 58272
rect 800 57992 119120 58128
rect 800 57592 119200 57992
rect 800 57456 119120 57592
rect 880 57312 119120 57456
rect 880 57176 119200 57312
rect 800 57048 119200 57176
rect 800 56768 119120 57048
rect 800 56504 119200 56768
rect 880 56368 119200 56504
rect 880 56224 119120 56368
rect 800 56088 119120 56224
rect 800 55688 119200 56088
rect 800 55552 119120 55688
rect 880 55408 119120 55552
rect 880 55272 119200 55408
rect 800 55144 119200 55272
rect 800 54864 119120 55144
rect 800 54600 119200 54864
rect 880 54464 119200 54600
rect 880 54320 119120 54464
rect 800 54184 119120 54320
rect 800 53920 119200 54184
rect 800 53648 119120 53920
rect 880 53640 119120 53648
rect 880 53368 119200 53640
rect 800 53240 119200 53368
rect 800 52960 119120 53240
rect 800 52696 119200 52960
rect 880 52560 119200 52696
rect 880 52416 119120 52560
rect 800 52280 119120 52416
rect 800 52016 119200 52280
rect 800 51744 119120 52016
rect 880 51736 119120 51744
rect 880 51464 119200 51736
rect 800 51336 119200 51464
rect 800 51056 119120 51336
rect 800 50792 119200 51056
rect 880 50512 119120 50792
rect 800 50112 119200 50512
rect 800 49840 119120 50112
rect 880 49832 119120 49840
rect 880 49560 119200 49832
rect 800 49432 119200 49560
rect 800 49152 119120 49432
rect 800 48888 119200 49152
rect 880 48608 119120 48888
rect 800 48208 119200 48608
rect 800 47936 119120 48208
rect 880 47928 119120 47936
rect 880 47664 119200 47928
rect 880 47656 119120 47664
rect 800 47384 119120 47656
rect 800 46984 119200 47384
rect 880 46704 119120 46984
rect 800 46304 119200 46704
rect 800 46032 119120 46304
rect 880 46024 119120 46032
rect 880 45760 119200 46024
rect 880 45752 119120 45760
rect 800 45480 119120 45752
rect 800 45080 119200 45480
rect 880 44800 119120 45080
rect 800 44536 119200 44800
rect 800 44256 119120 44536
rect 800 44128 119200 44256
rect 880 43856 119200 44128
rect 880 43848 119120 43856
rect 800 43576 119120 43848
rect 800 43176 119200 43576
rect 880 42896 119120 43176
rect 800 42632 119200 42896
rect 800 42352 119120 42632
rect 800 42224 119200 42352
rect 880 41952 119200 42224
rect 880 41944 119120 41952
rect 800 41672 119120 41944
rect 800 41408 119200 41672
rect 800 41272 119120 41408
rect 880 41128 119120 41272
rect 880 40992 119200 41128
rect 800 40728 119200 40992
rect 800 40448 119120 40728
rect 800 40320 119200 40448
rect 880 40184 119200 40320
rect 880 40040 119120 40184
rect 800 39904 119120 40040
rect 800 39504 119200 39904
rect 800 39368 119120 39504
rect 880 39224 119120 39368
rect 880 39088 119200 39224
rect 800 38824 119200 39088
rect 800 38544 119120 38824
rect 800 38416 119200 38544
rect 880 38280 119200 38416
rect 880 38136 119120 38280
rect 800 38000 119120 38136
rect 800 37600 119200 38000
rect 800 37464 119120 37600
rect 880 37320 119120 37464
rect 880 37184 119200 37320
rect 800 37056 119200 37184
rect 800 36776 119120 37056
rect 800 36512 119200 36776
rect 880 36376 119200 36512
rect 880 36232 119120 36376
rect 800 36096 119120 36232
rect 800 35696 119200 36096
rect 800 35560 119120 35696
rect 880 35416 119120 35560
rect 880 35280 119200 35416
rect 800 35152 119200 35280
rect 800 34872 119120 35152
rect 800 34608 119200 34872
rect 880 34472 119200 34608
rect 880 34328 119120 34472
rect 800 34192 119120 34328
rect 800 33928 119200 34192
rect 800 33656 119120 33928
rect 880 33648 119120 33656
rect 880 33376 119200 33648
rect 800 33248 119200 33376
rect 800 32968 119120 33248
rect 800 32704 119200 32968
rect 880 32568 119200 32704
rect 880 32424 119120 32568
rect 800 32288 119120 32424
rect 800 32024 119200 32288
rect 800 31752 119120 32024
rect 880 31744 119120 31752
rect 880 31472 119200 31744
rect 800 31344 119200 31472
rect 800 31064 119120 31344
rect 800 30800 119200 31064
rect 880 30520 119120 30800
rect 800 30120 119200 30520
rect 800 29848 119120 30120
rect 880 29840 119120 29848
rect 880 29568 119200 29840
rect 800 29440 119200 29568
rect 800 29160 119120 29440
rect 800 28896 119200 29160
rect 880 28616 119120 28896
rect 800 28216 119200 28616
rect 800 27944 119120 28216
rect 880 27936 119120 27944
rect 880 27672 119200 27936
rect 880 27664 119120 27672
rect 800 27392 119120 27664
rect 800 26992 119200 27392
rect 880 26712 119120 26992
rect 800 26312 119200 26712
rect 800 26040 119120 26312
rect 880 26032 119120 26040
rect 880 25768 119200 26032
rect 880 25760 119120 25768
rect 800 25488 119120 25760
rect 800 25088 119200 25488
rect 880 24808 119120 25088
rect 800 24544 119200 24808
rect 800 24264 119120 24544
rect 800 24136 119200 24264
rect 880 23864 119200 24136
rect 880 23856 119120 23864
rect 800 23584 119120 23856
rect 800 23184 119200 23584
rect 880 22904 119120 23184
rect 800 22640 119200 22904
rect 800 22360 119120 22640
rect 800 22232 119200 22360
rect 880 21960 119200 22232
rect 880 21952 119120 21960
rect 800 21680 119120 21952
rect 800 21416 119200 21680
rect 800 21280 119120 21416
rect 880 21136 119120 21280
rect 880 21000 119200 21136
rect 800 20736 119200 21000
rect 800 20456 119120 20736
rect 800 20328 119200 20456
rect 880 20192 119200 20328
rect 880 20048 119120 20192
rect 800 19912 119120 20048
rect 800 19512 119200 19912
rect 800 19376 119120 19512
rect 880 19232 119120 19376
rect 880 19096 119200 19232
rect 800 18832 119200 19096
rect 800 18552 119120 18832
rect 800 18424 119200 18552
rect 880 18288 119200 18424
rect 880 18144 119120 18288
rect 800 18008 119120 18144
rect 800 17608 119200 18008
rect 800 17472 119120 17608
rect 880 17328 119120 17472
rect 880 17192 119200 17328
rect 800 17064 119200 17192
rect 800 16784 119120 17064
rect 800 16520 119200 16784
rect 880 16384 119200 16520
rect 880 16240 119120 16384
rect 800 16104 119120 16240
rect 800 15704 119200 16104
rect 800 15568 119120 15704
rect 880 15424 119120 15568
rect 880 15288 119200 15424
rect 800 15160 119200 15288
rect 800 14880 119120 15160
rect 800 14616 119200 14880
rect 880 14480 119200 14616
rect 880 14336 119120 14480
rect 800 14200 119120 14336
rect 800 13936 119200 14200
rect 800 13664 119120 13936
rect 880 13656 119120 13664
rect 880 13384 119200 13656
rect 800 13256 119200 13384
rect 800 12976 119120 13256
rect 800 12712 119200 12976
rect 880 12576 119200 12712
rect 880 12432 119120 12576
rect 800 12296 119120 12432
rect 800 12032 119200 12296
rect 800 11760 119120 12032
rect 880 11752 119120 11760
rect 880 11480 119200 11752
rect 800 11352 119200 11480
rect 800 11072 119120 11352
rect 800 10808 119200 11072
rect 880 10528 119120 10808
rect 800 10128 119200 10528
rect 800 9856 119120 10128
rect 880 9848 119120 9856
rect 880 9576 119200 9848
rect 800 9448 119200 9576
rect 800 9168 119120 9448
rect 800 8904 119200 9168
rect 880 8624 119120 8904
rect 800 8224 119200 8624
rect 800 7952 119120 8224
rect 880 7944 119120 7952
rect 880 7680 119200 7944
rect 880 7672 119120 7680
rect 800 7400 119120 7672
rect 800 7000 119200 7400
rect 880 6720 119120 7000
rect 800 6320 119200 6720
rect 800 6048 119120 6320
rect 880 6040 119120 6048
rect 880 5776 119200 6040
rect 880 5768 119120 5776
rect 800 5496 119120 5768
rect 800 5096 119200 5496
rect 880 4816 119120 5096
rect 800 4552 119200 4816
rect 800 4272 119120 4552
rect 800 4144 119200 4272
rect 880 3872 119200 4144
rect 880 3864 119120 3872
rect 800 3592 119120 3864
rect 800 3192 119200 3592
rect 880 2912 119120 3192
rect 800 2648 119200 2912
rect 800 2368 119120 2648
rect 800 2240 119200 2368
rect 880 1968 119200 2240
rect 880 1960 119120 1968
rect 800 1688 119120 1960
rect 800 1424 119200 1688
rect 800 1288 119120 1424
rect 880 1144 119120 1288
rect 880 1008 119200 1144
rect 800 744 119200 1008
rect 800 464 119120 744
rect 800 336 119200 464
rect 880 200 119200 336
rect 880 56 119120 200
rect 800 27 119120 56
<< metal4 >>
rect 4208 1848 4528 77560
rect 19568 1848 19888 77560
rect 34928 1848 35248 77560
rect 50288 1848 50608 77560
rect 65648 1848 65968 77560
rect 81008 1848 81328 77560
rect 96368 1848 96688 77560
rect 111728 1848 112048 77560
<< obsm4 >>
rect 2819 3291 4128 76117
rect 4608 3291 19488 76117
rect 19968 3291 34848 76117
rect 35328 3291 50208 76117
rect 50688 3291 65568 76117
rect 66048 3291 80928 76117
rect 81408 3291 96288 76117
rect 96768 3291 111648 76117
rect 112128 3291 116045 76117
<< labels >>
rlabel metal3 s 0 3944 800 4064 6 A[0]
port 1 nsew signal input
rlabel metal3 s 0 13464 800 13584 6 A[10]
port 2 nsew signal input
rlabel metal3 s 0 14416 800 14536 6 A[11]
port 3 nsew signal input
rlabel metal3 s 0 15368 800 15488 6 A[12]
port 4 nsew signal input
rlabel metal3 s 0 16320 800 16440 6 A[13]
port 5 nsew signal input
rlabel metal3 s 0 17272 800 17392 6 A[14]
port 6 nsew signal input
rlabel metal3 s 0 18224 800 18344 6 A[15]
port 7 nsew signal input
rlabel metal3 s 0 19176 800 19296 6 A[16]
port 8 nsew signal input
rlabel metal3 s 0 20128 800 20248 6 A[17]
port 9 nsew signal input
rlabel metal3 s 0 21080 800 21200 6 A[18]
port 10 nsew signal input
rlabel metal3 s 0 22032 800 22152 6 A[19]
port 11 nsew signal input
rlabel metal3 s 0 4896 800 5016 6 A[1]
port 12 nsew signal input
rlabel metal3 s 0 22984 800 23104 6 A[20]
port 13 nsew signal input
rlabel metal3 s 0 23936 800 24056 6 A[21]
port 14 nsew signal input
rlabel metal3 s 0 24888 800 25008 6 A[22]
port 15 nsew signal input
rlabel metal3 s 0 25840 800 25960 6 A[23]
port 16 nsew signal input
rlabel metal3 s 0 5848 800 5968 6 A[2]
port 17 nsew signal input
rlabel metal3 s 0 6800 800 6920 6 A[3]
port 18 nsew signal input
rlabel metal3 s 0 7752 800 7872 6 A[4]
port 19 nsew signal input
rlabel metal3 s 0 8704 800 8824 6 A[5]
port 20 nsew signal input
rlabel metal3 s 0 9656 800 9776 6 A[6]
port 21 nsew signal input
rlabel metal3 s 0 10608 800 10728 6 A[7]
port 22 nsew signal input
rlabel metal3 s 0 11560 800 11680 6 A[8]
port 23 nsew signal input
rlabel metal3 s 0 12512 800 12632 6 A[9]
port 24 nsew signal input
rlabel metal3 s 0 26792 800 26912 6 A_h[0]
port 25 nsew signal input
rlabel metal3 s 0 36312 800 36432 6 A_h[10]
port 26 nsew signal input
rlabel metal3 s 0 37264 800 37384 6 A_h[11]
port 27 nsew signal input
rlabel metal3 s 0 38216 800 38336 6 A_h[12]
port 28 nsew signal input
rlabel metal3 s 0 39168 800 39288 6 A_h[13]
port 29 nsew signal input
rlabel metal3 s 0 40120 800 40240 6 A_h[14]
port 30 nsew signal input
rlabel metal3 s 0 41072 800 41192 6 A_h[15]
port 31 nsew signal input
rlabel metal3 s 0 42024 800 42144 6 A_h[16]
port 32 nsew signal input
rlabel metal3 s 0 42976 800 43096 6 A_h[17]
port 33 nsew signal input
rlabel metal3 s 0 43928 800 44048 6 A_h[18]
port 34 nsew signal input
rlabel metal3 s 0 44880 800 45000 6 A_h[19]
port 35 nsew signal input
rlabel metal3 s 0 27744 800 27864 6 A_h[1]
port 36 nsew signal input
rlabel metal3 s 0 45832 800 45952 6 A_h[20]
port 37 nsew signal input
rlabel metal3 s 0 46784 800 46904 6 A_h[21]
port 38 nsew signal input
rlabel metal3 s 0 47736 800 47856 6 A_h[22]
port 39 nsew signal input
rlabel metal3 s 0 48688 800 48808 6 A_h[23]
port 40 nsew signal input
rlabel metal3 s 0 28696 800 28816 6 A_h[2]
port 41 nsew signal input
rlabel metal3 s 0 29648 800 29768 6 A_h[3]
port 42 nsew signal input
rlabel metal3 s 0 30600 800 30720 6 A_h[4]
port 43 nsew signal input
rlabel metal3 s 0 31552 800 31672 6 A_h[5]
port 44 nsew signal input
rlabel metal3 s 0 32504 800 32624 6 A_h[6]
port 45 nsew signal input
rlabel metal3 s 0 33456 800 33576 6 A_h[7]
port 46 nsew signal input
rlabel metal3 s 0 34408 800 34528 6 A_h[8]
port 47 nsew signal input
rlabel metal3 s 0 35360 800 35480 6 A_h[9]
port 48 nsew signal input
rlabel metal3 s 0 49640 800 49760 6 Do[0]
port 49 nsew signal output
rlabel metal3 s 0 59160 800 59280 6 Do[10]
port 50 nsew signal output
rlabel metal3 s 0 60112 800 60232 6 Do[11]
port 51 nsew signal output
rlabel metal3 s 0 61064 800 61184 6 Do[12]
port 52 nsew signal output
rlabel metal3 s 0 62016 800 62136 6 Do[13]
port 53 nsew signal output
rlabel metal3 s 0 62968 800 63088 6 Do[14]
port 54 nsew signal output
rlabel metal3 s 0 63920 800 64040 6 Do[15]
port 55 nsew signal output
rlabel metal3 s 0 64872 800 64992 6 Do[16]
port 56 nsew signal output
rlabel metal3 s 0 65824 800 65944 6 Do[17]
port 57 nsew signal output
rlabel metal3 s 0 66776 800 66896 6 Do[18]
port 58 nsew signal output
rlabel metal3 s 0 67728 800 67848 6 Do[19]
port 59 nsew signal output
rlabel metal3 s 0 50592 800 50712 6 Do[1]
port 60 nsew signal output
rlabel metal3 s 0 68680 800 68800 6 Do[20]
port 61 nsew signal output
rlabel metal3 s 0 69632 800 69752 6 Do[21]
port 62 nsew signal output
rlabel metal3 s 0 70584 800 70704 6 Do[22]
port 63 nsew signal output
rlabel metal3 s 0 71536 800 71656 6 Do[23]
port 64 nsew signal output
rlabel metal3 s 0 72488 800 72608 6 Do[24]
port 65 nsew signal output
rlabel metal3 s 0 73440 800 73560 6 Do[25]
port 66 nsew signal output
rlabel metal3 s 0 74392 800 74512 6 Do[26]
port 67 nsew signal output
rlabel metal3 s 0 75344 800 75464 6 Do[27]
port 68 nsew signal output
rlabel metal3 s 0 76296 800 76416 6 Do[28]
port 69 nsew signal output
rlabel metal3 s 0 77248 800 77368 6 Do[29]
port 70 nsew signal output
rlabel metal3 s 0 51544 800 51664 6 Do[2]
port 71 nsew signal output
rlabel metal3 s 0 78200 800 78320 6 Do[30]
port 72 nsew signal output
rlabel metal3 s 0 79152 800 79272 6 Do[31]
port 73 nsew signal output
rlabel metal3 s 0 52496 800 52616 6 Do[3]
port 74 nsew signal output
rlabel metal3 s 0 53448 800 53568 6 Do[4]
port 75 nsew signal output
rlabel metal3 s 0 54400 800 54520 6 Do[5]
port 76 nsew signal output
rlabel metal3 s 0 55352 800 55472 6 Do[6]
port 77 nsew signal output
rlabel metal3 s 0 56304 800 56424 6 Do[7]
port 78 nsew signal output
rlabel metal3 s 0 57256 800 57376 6 Do[8]
port 79 nsew signal output
rlabel metal3 s 0 58208 800 58328 6 Do[9]
port 80 nsew signal output
rlabel metal3 s 0 136 800 256 6 clk
port 81 nsew signal input
rlabel metal3 s 0 2992 800 3112 6 hit
port 82 nsew signal output
rlabel metal3 s 119200 0 120000 120 6 line[0]
port 83 nsew signal input
rlabel metal3 s 119200 62424 120000 62544 6 line[100]
port 84 nsew signal input
rlabel metal3 s 119200 62968 120000 63088 6 line[101]
port 85 nsew signal input
rlabel metal3 s 119200 63648 120000 63768 6 line[102]
port 86 nsew signal input
rlabel metal3 s 119200 64328 120000 64448 6 line[103]
port 87 nsew signal input
rlabel metal3 s 119200 64872 120000 64992 6 line[104]
port 88 nsew signal input
rlabel metal3 s 119200 65552 120000 65672 6 line[105]
port 89 nsew signal input
rlabel metal3 s 119200 66096 120000 66216 6 line[106]
port 90 nsew signal input
rlabel metal3 s 119200 66776 120000 66896 6 line[107]
port 91 nsew signal input
rlabel metal3 s 119200 67456 120000 67576 6 line[108]
port 92 nsew signal input
rlabel metal3 s 119200 68000 120000 68120 6 line[109]
port 93 nsew signal input
rlabel metal3 s 119200 6120 120000 6240 6 line[10]
port 94 nsew signal input
rlabel metal3 s 119200 68680 120000 68800 6 line[110]
port 95 nsew signal input
rlabel metal3 s 119200 69224 120000 69344 6 line[111]
port 96 nsew signal input
rlabel metal3 s 119200 69904 120000 70024 6 line[112]
port 97 nsew signal input
rlabel metal3 s 119200 70584 120000 70704 6 line[113]
port 98 nsew signal input
rlabel metal3 s 119200 71128 120000 71248 6 line[114]
port 99 nsew signal input
rlabel metal3 s 119200 71808 120000 71928 6 line[115]
port 100 nsew signal input
rlabel metal3 s 119200 72352 120000 72472 6 line[116]
port 101 nsew signal input
rlabel metal3 s 119200 73032 120000 73152 6 line[117]
port 102 nsew signal input
rlabel metal3 s 119200 73712 120000 73832 6 line[118]
port 103 nsew signal input
rlabel metal3 s 119200 74256 120000 74376 6 line[119]
port 104 nsew signal input
rlabel metal3 s 119200 6800 120000 6920 6 line[11]
port 105 nsew signal input
rlabel metal3 s 119200 74936 120000 75056 6 line[120]
port 106 nsew signal input
rlabel metal3 s 119200 75480 120000 75600 6 line[121]
port 107 nsew signal input
rlabel metal3 s 119200 76160 120000 76280 6 line[122]
port 108 nsew signal input
rlabel metal3 s 119200 76840 120000 76960 6 line[123]
port 109 nsew signal input
rlabel metal3 s 119200 77384 120000 77504 6 line[124]
port 110 nsew signal input
rlabel metal3 s 119200 78064 120000 78184 6 line[125]
port 111 nsew signal input
rlabel metal3 s 119200 78608 120000 78728 6 line[126]
port 112 nsew signal input
rlabel metal3 s 119200 79288 120000 79408 6 line[127]
port 113 nsew signal input
rlabel metal3 s 119200 7480 120000 7600 6 line[12]
port 114 nsew signal input
rlabel metal3 s 119200 8024 120000 8144 6 line[13]
port 115 nsew signal input
rlabel metal3 s 119200 8704 120000 8824 6 line[14]
port 116 nsew signal input
rlabel metal3 s 119200 9248 120000 9368 6 line[15]
port 117 nsew signal input
rlabel metal3 s 119200 9928 120000 10048 6 line[16]
port 118 nsew signal input
rlabel metal3 s 119200 10608 120000 10728 6 line[17]
port 119 nsew signal input
rlabel metal3 s 119200 11152 120000 11272 6 line[18]
port 120 nsew signal input
rlabel metal3 s 119200 11832 120000 11952 6 line[19]
port 121 nsew signal input
rlabel metal3 s 119200 544 120000 664 6 line[1]
port 122 nsew signal input
rlabel metal3 s 119200 12376 120000 12496 6 line[20]
port 123 nsew signal input
rlabel metal3 s 119200 13056 120000 13176 6 line[21]
port 124 nsew signal input
rlabel metal3 s 119200 13736 120000 13856 6 line[22]
port 125 nsew signal input
rlabel metal3 s 119200 14280 120000 14400 6 line[23]
port 126 nsew signal input
rlabel metal3 s 119200 14960 120000 15080 6 line[24]
port 127 nsew signal input
rlabel metal3 s 119200 15504 120000 15624 6 line[25]
port 128 nsew signal input
rlabel metal3 s 119200 16184 120000 16304 6 line[26]
port 129 nsew signal input
rlabel metal3 s 119200 16864 120000 16984 6 line[27]
port 130 nsew signal input
rlabel metal3 s 119200 17408 120000 17528 6 line[28]
port 131 nsew signal input
rlabel metal3 s 119200 18088 120000 18208 6 line[29]
port 132 nsew signal input
rlabel metal3 s 119200 1224 120000 1344 6 line[2]
port 133 nsew signal input
rlabel metal3 s 119200 18632 120000 18752 6 line[30]
port 134 nsew signal input
rlabel metal3 s 119200 19312 120000 19432 6 line[31]
port 135 nsew signal input
rlabel metal3 s 119200 19992 120000 20112 6 line[32]
port 136 nsew signal input
rlabel metal3 s 119200 20536 120000 20656 6 line[33]
port 137 nsew signal input
rlabel metal3 s 119200 21216 120000 21336 6 line[34]
port 138 nsew signal input
rlabel metal3 s 119200 21760 120000 21880 6 line[35]
port 139 nsew signal input
rlabel metal3 s 119200 22440 120000 22560 6 line[36]
port 140 nsew signal input
rlabel metal3 s 119200 22984 120000 23104 6 line[37]
port 141 nsew signal input
rlabel metal3 s 119200 23664 120000 23784 6 line[38]
port 142 nsew signal input
rlabel metal3 s 119200 24344 120000 24464 6 line[39]
port 143 nsew signal input
rlabel metal3 s 119200 1768 120000 1888 6 line[3]
port 144 nsew signal input
rlabel metal3 s 119200 24888 120000 25008 6 line[40]
port 145 nsew signal input
rlabel metal3 s 119200 25568 120000 25688 6 line[41]
port 146 nsew signal input
rlabel metal3 s 119200 26112 120000 26232 6 line[42]
port 147 nsew signal input
rlabel metal3 s 119200 26792 120000 26912 6 line[43]
port 148 nsew signal input
rlabel metal3 s 119200 27472 120000 27592 6 line[44]
port 149 nsew signal input
rlabel metal3 s 119200 28016 120000 28136 6 line[45]
port 150 nsew signal input
rlabel metal3 s 119200 28696 120000 28816 6 line[46]
port 151 nsew signal input
rlabel metal3 s 119200 29240 120000 29360 6 line[47]
port 152 nsew signal input
rlabel metal3 s 119200 29920 120000 30040 6 line[48]
port 153 nsew signal input
rlabel metal3 s 119200 30600 120000 30720 6 line[49]
port 154 nsew signal input
rlabel metal3 s 119200 2448 120000 2568 6 line[4]
port 155 nsew signal input
rlabel metal3 s 119200 31144 120000 31264 6 line[50]
port 156 nsew signal input
rlabel metal3 s 119200 31824 120000 31944 6 line[51]
port 157 nsew signal input
rlabel metal3 s 119200 32368 120000 32488 6 line[52]
port 158 nsew signal input
rlabel metal3 s 119200 33048 120000 33168 6 line[53]
port 159 nsew signal input
rlabel metal3 s 119200 33728 120000 33848 6 line[54]
port 160 nsew signal input
rlabel metal3 s 119200 34272 120000 34392 6 line[55]
port 161 nsew signal input
rlabel metal3 s 119200 34952 120000 35072 6 line[56]
port 162 nsew signal input
rlabel metal3 s 119200 35496 120000 35616 6 line[57]
port 163 nsew signal input
rlabel metal3 s 119200 36176 120000 36296 6 line[58]
port 164 nsew signal input
rlabel metal3 s 119200 36856 120000 36976 6 line[59]
port 165 nsew signal input
rlabel metal3 s 119200 2992 120000 3112 6 line[5]
port 166 nsew signal input
rlabel metal3 s 119200 37400 120000 37520 6 line[60]
port 167 nsew signal input
rlabel metal3 s 119200 38080 120000 38200 6 line[61]
port 168 nsew signal input
rlabel metal3 s 119200 38624 120000 38744 6 line[62]
port 169 nsew signal input
rlabel metal3 s 119200 39304 120000 39424 6 line[63]
port 170 nsew signal input
rlabel metal3 s 119200 39984 120000 40104 6 line[64]
port 171 nsew signal input
rlabel metal3 s 119200 40528 120000 40648 6 line[65]
port 172 nsew signal input
rlabel metal3 s 119200 41208 120000 41328 6 line[66]
port 173 nsew signal input
rlabel metal3 s 119200 41752 120000 41872 6 line[67]
port 174 nsew signal input
rlabel metal3 s 119200 42432 120000 42552 6 line[68]
port 175 nsew signal input
rlabel metal3 s 119200 42976 120000 43096 6 line[69]
port 176 nsew signal input
rlabel metal3 s 119200 3672 120000 3792 6 line[6]
port 177 nsew signal input
rlabel metal3 s 119200 43656 120000 43776 6 line[70]
port 178 nsew signal input
rlabel metal3 s 119200 44336 120000 44456 6 line[71]
port 179 nsew signal input
rlabel metal3 s 119200 44880 120000 45000 6 line[72]
port 180 nsew signal input
rlabel metal3 s 119200 45560 120000 45680 6 line[73]
port 181 nsew signal input
rlabel metal3 s 119200 46104 120000 46224 6 line[74]
port 182 nsew signal input
rlabel metal3 s 119200 46784 120000 46904 6 line[75]
port 183 nsew signal input
rlabel metal3 s 119200 47464 120000 47584 6 line[76]
port 184 nsew signal input
rlabel metal3 s 119200 48008 120000 48128 6 line[77]
port 185 nsew signal input
rlabel metal3 s 119200 48688 120000 48808 6 line[78]
port 186 nsew signal input
rlabel metal3 s 119200 49232 120000 49352 6 line[79]
port 187 nsew signal input
rlabel metal3 s 119200 4352 120000 4472 6 line[7]
port 188 nsew signal input
rlabel metal3 s 119200 49912 120000 50032 6 line[80]
port 189 nsew signal input
rlabel metal3 s 119200 50592 120000 50712 6 line[81]
port 190 nsew signal input
rlabel metal3 s 119200 51136 120000 51256 6 line[82]
port 191 nsew signal input
rlabel metal3 s 119200 51816 120000 51936 6 line[83]
port 192 nsew signal input
rlabel metal3 s 119200 52360 120000 52480 6 line[84]
port 193 nsew signal input
rlabel metal3 s 119200 53040 120000 53160 6 line[85]
port 194 nsew signal input
rlabel metal3 s 119200 53720 120000 53840 6 line[86]
port 195 nsew signal input
rlabel metal3 s 119200 54264 120000 54384 6 line[87]
port 196 nsew signal input
rlabel metal3 s 119200 54944 120000 55064 6 line[88]
port 197 nsew signal input
rlabel metal3 s 119200 55488 120000 55608 6 line[89]
port 198 nsew signal input
rlabel metal3 s 119200 4896 120000 5016 6 line[8]
port 199 nsew signal input
rlabel metal3 s 119200 56168 120000 56288 6 line[90]
port 200 nsew signal input
rlabel metal3 s 119200 56848 120000 56968 6 line[91]
port 201 nsew signal input
rlabel metal3 s 119200 57392 120000 57512 6 line[92]
port 202 nsew signal input
rlabel metal3 s 119200 58072 120000 58192 6 line[93]
port 203 nsew signal input
rlabel metal3 s 119200 58616 120000 58736 6 line[94]
port 204 nsew signal input
rlabel metal3 s 119200 59296 120000 59416 6 line[95]
port 205 nsew signal input
rlabel metal3 s 119200 59976 120000 60096 6 line[96]
port 206 nsew signal input
rlabel metal3 s 119200 60520 120000 60640 6 line[97]
port 207 nsew signal input
rlabel metal3 s 119200 61200 120000 61320 6 line[98]
port 208 nsew signal input
rlabel metal3 s 119200 61744 120000 61864 6 line[99]
port 209 nsew signal input
rlabel metal3 s 119200 5576 120000 5696 6 line[9]
port 210 nsew signal input
rlabel metal3 s 0 1088 800 1208 6 rst_n
port 211 nsew signal input
rlabel metal3 s 0 2040 800 2160 6 wr
port 212 nsew signal input
rlabel metal4 s 96368 1848 96688 77560 6 VPWR
port 213 nsew power bidirectional
rlabel metal4 s 65648 1848 65968 77560 6 VPWR
port 214 nsew power bidirectional
rlabel metal4 s 34928 1848 35248 77560 6 VPWR
port 215 nsew power bidirectional
rlabel metal4 s 4208 1848 4528 77560 6 VPWR
port 216 nsew power bidirectional
rlabel metal4 s 111728 1848 112048 77560 6 VGND
port 217 nsew ground bidirectional
rlabel metal4 s 81008 1848 81328 77560 6 VGND
port 218 nsew ground bidirectional
rlabel metal4 s 50288 1848 50608 77560 6 VGND
port 219 nsew ground bidirectional
rlabel metal4 s 19568 1848 19888 77560 6 VGND
port 220 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 120000 79408
string LEFview TRUE
<< end >>
