VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DMC_32x16HC
  CLASS BLOCK ;
  FOREIGN DMC_32x16HC ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 397.040 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.720 4.000 20.320 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.320 4.000 67.920 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.080 4.000 72.680 ;
    END
  END A[11]
  PIN A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.840 4.000 77.440 ;
    END
  END A[12]
  PIN A[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.600 4.000 82.200 ;
    END
  END A[13]
  PIN A[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.360 4.000 86.960 ;
    END
  END A[14]
  PIN A[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.120 4.000 91.720 ;
    END
  END A[15]
  PIN A[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.880 4.000 96.480 ;
    END
  END A[16]
  PIN A[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.640 4.000 101.240 ;
    END
  END A[17]
  PIN A[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.400 4.000 106.000 ;
    END
  END A[18]
  PIN A[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.160 4.000 110.760 ;
    END
  END A[19]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.480 4.000 25.080 ;
    END
  END A[1]
  PIN A[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.920 4.000 115.520 ;
    END
  END A[20]
  PIN A[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.680 4.000 120.280 ;
    END
  END A[21]
  PIN A[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.440 4.000 125.040 ;
    END
  END A[22]
  PIN A[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.200 4.000 129.800 ;
    END
  END A[23]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.240 4.000 29.840 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.000 4.000 34.600 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.760 4.000 39.360 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.520 4.000 44.120 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.280 4.000 48.880 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.040 4.000 53.640 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.800 4.000 58.400 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.560 4.000 63.160 ;
    END
  END A[9]
  PIN A_h[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.960 4.000 134.560 ;
    END
  END A_h[0]
  PIN A_h[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.560 4.000 182.160 ;
    END
  END A_h[10]
  PIN A_h[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.320 4.000 186.920 ;
    END
  END A_h[11]
  PIN A_h[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.080 4.000 191.680 ;
    END
  END A_h[12]
  PIN A_h[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.840 4.000 196.440 ;
    END
  END A_h[13]
  PIN A_h[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.600 4.000 201.200 ;
    END
  END A_h[14]
  PIN A_h[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.360 4.000 205.960 ;
    END
  END A_h[15]
  PIN A_h[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.120 4.000 210.720 ;
    END
  END A_h[16]
  PIN A_h[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.880 4.000 215.480 ;
    END
  END A_h[17]
  PIN A_h[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.640 4.000 220.240 ;
    END
  END A_h[18]
  PIN A_h[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.400 4.000 225.000 ;
    END
  END A_h[19]
  PIN A_h[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.720 4.000 139.320 ;
    END
  END A_h[1]
  PIN A_h[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.160 4.000 229.760 ;
    END
  END A_h[20]
  PIN A_h[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.920 4.000 234.520 ;
    END
  END A_h[21]
  PIN A_h[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.680 4.000 239.280 ;
    END
  END A_h[22]
  PIN A_h[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.440 4.000 244.040 ;
    END
  END A_h[23]
  PIN A_h[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.480 4.000 144.080 ;
    END
  END A_h[2]
  PIN A_h[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.240 4.000 148.840 ;
    END
  END A_h[3]
  PIN A_h[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.000 4.000 153.600 ;
    END
  END A_h[4]
  PIN A_h[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.760 4.000 158.360 ;
    END
  END A_h[5]
  PIN A_h[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.520 4.000 163.120 ;
    END
  END A_h[6]
  PIN A_h[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.280 4.000 167.880 ;
    END
  END A_h[7]
  PIN A_h[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.040 4.000 172.640 ;
    END
  END A_h[8]
  PIN A_h[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.800 4.000 177.400 ;
    END
  END A_h[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.200 4.000 248.800 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.800 4.000 296.400 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.560 4.000 301.160 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.320 4.000 305.920 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.080 4.000 310.680 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.840 4.000 315.440 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.600 4.000 320.200 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.360 4.000 324.960 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.120 4.000 329.720 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.880 4.000 334.480 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.640 4.000 339.240 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.960 4.000 253.560 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.400 4.000 344.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.160 4.000 348.760 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.920 4.000 353.520 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.680 4.000 358.280 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.440 4.000 363.040 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.200 4.000 367.800 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.960 4.000 372.560 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.720 4.000 377.320 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.480 4.000 382.080 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.240 4.000 386.840 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.720 4.000 258.320 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.000 4.000 391.600 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.760 4.000 396.360 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.480 4.000 263.080 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.240 4.000 267.840 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.000 4.000 272.600 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.760 4.000 277.360 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.520 4.000 282.120 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.280 4.000 286.880 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.040 4.000 291.640 ;
    END
  END Do[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.680 4.000 1.280 ;
    END
  END clk
  PIN hit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.960 4.000 15.560 ;
    END
  END hit
  PIN line[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 0.000 600.000 0.600 ;
    END
  END line[0]
  PIN line[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 312.120 600.000 312.720 ;
    END
  END line[100]
  PIN line[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 314.840 600.000 315.440 ;
    END
  END line[101]
  PIN line[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 318.240 600.000 318.840 ;
    END
  END line[102]
  PIN line[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 321.640 600.000 322.240 ;
    END
  END line[103]
  PIN line[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 324.360 600.000 324.960 ;
    END
  END line[104]
  PIN line[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 327.760 600.000 328.360 ;
    END
  END line[105]
  PIN line[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 330.480 600.000 331.080 ;
    END
  END line[106]
  PIN line[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 333.880 600.000 334.480 ;
    END
  END line[107]
  PIN line[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 337.280 600.000 337.880 ;
    END
  END line[108]
  PIN line[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 340.000 600.000 340.600 ;
    END
  END line[109]
  PIN line[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 30.600 600.000 31.200 ;
    END
  END line[10]
  PIN line[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 343.400 600.000 344.000 ;
    END
  END line[110]
  PIN line[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 346.120 600.000 346.720 ;
    END
  END line[111]
  PIN line[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 349.520 600.000 350.120 ;
    END
  END line[112]
  PIN line[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 352.920 600.000 353.520 ;
    END
  END line[113]
  PIN line[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 355.640 600.000 356.240 ;
    END
  END line[114]
  PIN line[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 359.040 600.000 359.640 ;
    END
  END line[115]
  PIN line[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 361.760 600.000 362.360 ;
    END
  END line[116]
  PIN line[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 365.160 600.000 365.760 ;
    END
  END line[117]
  PIN line[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 368.560 600.000 369.160 ;
    END
  END line[118]
  PIN line[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 371.280 600.000 371.880 ;
    END
  END line[119]
  PIN line[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 34.000 600.000 34.600 ;
    END
  END line[11]
  PIN line[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 374.680 600.000 375.280 ;
    END
  END line[120]
  PIN line[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 377.400 600.000 378.000 ;
    END
  END line[121]
  PIN line[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 380.800 600.000 381.400 ;
    END
  END line[122]
  PIN line[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 384.200 600.000 384.800 ;
    END
  END line[123]
  PIN line[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 386.920 600.000 387.520 ;
    END
  END line[124]
  PIN line[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 390.320 600.000 390.920 ;
    END
  END line[125]
  PIN line[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 393.040 600.000 393.640 ;
    END
  END line[126]
  PIN line[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 396.440 600.000 397.040 ;
    END
  END line[127]
  PIN line[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 37.400 600.000 38.000 ;
    END
  END line[12]
  PIN line[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 40.120 600.000 40.720 ;
    END
  END line[13]
  PIN line[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 43.520 600.000 44.120 ;
    END
  END line[14]
  PIN line[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 46.240 600.000 46.840 ;
    END
  END line[15]
  PIN line[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 49.640 600.000 50.240 ;
    END
  END line[16]
  PIN line[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 53.040 600.000 53.640 ;
    END
  END line[17]
  PIN line[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 55.760 600.000 56.360 ;
    END
  END line[18]
  PIN line[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 59.160 600.000 59.760 ;
    END
  END line[19]
  PIN line[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 2.720 600.000 3.320 ;
    END
  END line[1]
  PIN line[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 61.880 600.000 62.480 ;
    END
  END line[20]
  PIN line[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 65.280 600.000 65.880 ;
    END
  END line[21]
  PIN line[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 68.680 600.000 69.280 ;
    END
  END line[22]
  PIN line[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 71.400 600.000 72.000 ;
    END
  END line[23]
  PIN line[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 74.800 600.000 75.400 ;
    END
  END line[24]
  PIN line[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 77.520 600.000 78.120 ;
    END
  END line[25]
  PIN line[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 80.920 600.000 81.520 ;
    END
  END line[26]
  PIN line[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 84.320 600.000 84.920 ;
    END
  END line[27]
  PIN line[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 87.040 600.000 87.640 ;
    END
  END line[28]
  PIN line[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 90.440 600.000 91.040 ;
    END
  END line[29]
  PIN line[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 6.120 600.000 6.720 ;
    END
  END line[2]
  PIN line[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 93.160 600.000 93.760 ;
    END
  END line[30]
  PIN line[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 96.560 600.000 97.160 ;
    END
  END line[31]
  PIN line[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 99.960 600.000 100.560 ;
    END
  END line[32]
  PIN line[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 102.680 600.000 103.280 ;
    END
  END line[33]
  PIN line[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 106.080 600.000 106.680 ;
    END
  END line[34]
  PIN line[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 108.800 600.000 109.400 ;
    END
  END line[35]
  PIN line[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 112.200 600.000 112.800 ;
    END
  END line[36]
  PIN line[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 114.920 600.000 115.520 ;
    END
  END line[37]
  PIN line[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 118.320 600.000 118.920 ;
    END
  END line[38]
  PIN line[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 121.720 600.000 122.320 ;
    END
  END line[39]
  PIN line[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 8.840 600.000 9.440 ;
    END
  END line[3]
  PIN line[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 124.440 600.000 125.040 ;
    END
  END line[40]
  PIN line[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 127.840 600.000 128.440 ;
    END
  END line[41]
  PIN line[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 130.560 600.000 131.160 ;
    END
  END line[42]
  PIN line[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 133.960 600.000 134.560 ;
    END
  END line[43]
  PIN line[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 137.360 600.000 137.960 ;
    END
  END line[44]
  PIN line[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 140.080 600.000 140.680 ;
    END
  END line[45]
  PIN line[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 143.480 600.000 144.080 ;
    END
  END line[46]
  PIN line[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 146.200 600.000 146.800 ;
    END
  END line[47]
  PIN line[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 149.600 600.000 150.200 ;
    END
  END line[48]
  PIN line[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 153.000 600.000 153.600 ;
    END
  END line[49]
  PIN line[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 12.240 600.000 12.840 ;
    END
  END line[4]
  PIN line[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 155.720 600.000 156.320 ;
    END
  END line[50]
  PIN line[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 159.120 600.000 159.720 ;
    END
  END line[51]
  PIN line[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 161.840 600.000 162.440 ;
    END
  END line[52]
  PIN line[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 165.240 600.000 165.840 ;
    END
  END line[53]
  PIN line[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 168.640 600.000 169.240 ;
    END
  END line[54]
  PIN line[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 171.360 600.000 171.960 ;
    END
  END line[55]
  PIN line[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 174.760 600.000 175.360 ;
    END
  END line[56]
  PIN line[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 177.480 600.000 178.080 ;
    END
  END line[57]
  PIN line[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 180.880 600.000 181.480 ;
    END
  END line[58]
  PIN line[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 184.280 600.000 184.880 ;
    END
  END line[59]
  PIN line[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 14.960 600.000 15.560 ;
    END
  END line[5]
  PIN line[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 187.000 600.000 187.600 ;
    END
  END line[60]
  PIN line[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 190.400 600.000 191.000 ;
    END
  END line[61]
  PIN line[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 193.120 600.000 193.720 ;
    END
  END line[62]
  PIN line[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 196.520 600.000 197.120 ;
    END
  END line[63]
  PIN line[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 199.920 600.000 200.520 ;
    END
  END line[64]
  PIN line[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 202.640 600.000 203.240 ;
    END
  END line[65]
  PIN line[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 206.040 600.000 206.640 ;
    END
  END line[66]
  PIN line[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 208.760 600.000 209.360 ;
    END
  END line[67]
  PIN line[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 212.160 600.000 212.760 ;
    END
  END line[68]
  PIN line[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 214.880 600.000 215.480 ;
    END
  END line[69]
  PIN line[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 18.360 600.000 18.960 ;
    END
  END line[6]
  PIN line[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 218.280 600.000 218.880 ;
    END
  END line[70]
  PIN line[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 221.680 600.000 222.280 ;
    END
  END line[71]
  PIN line[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 224.400 600.000 225.000 ;
    END
  END line[72]
  PIN line[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 227.800 600.000 228.400 ;
    END
  END line[73]
  PIN line[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 230.520 600.000 231.120 ;
    END
  END line[74]
  PIN line[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 233.920 600.000 234.520 ;
    END
  END line[75]
  PIN line[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 237.320 600.000 237.920 ;
    END
  END line[76]
  PIN line[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 240.040 600.000 240.640 ;
    END
  END line[77]
  PIN line[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 243.440 600.000 244.040 ;
    END
  END line[78]
  PIN line[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 246.160 600.000 246.760 ;
    END
  END line[79]
  PIN line[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 21.760 600.000 22.360 ;
    END
  END line[7]
  PIN line[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 249.560 600.000 250.160 ;
    END
  END line[80]
  PIN line[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 252.960 600.000 253.560 ;
    END
  END line[81]
  PIN line[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 255.680 600.000 256.280 ;
    END
  END line[82]
  PIN line[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 259.080 600.000 259.680 ;
    END
  END line[83]
  PIN line[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 261.800 600.000 262.400 ;
    END
  END line[84]
  PIN line[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 265.200 600.000 265.800 ;
    END
  END line[85]
  PIN line[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 268.600 600.000 269.200 ;
    END
  END line[86]
  PIN line[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 271.320 600.000 271.920 ;
    END
  END line[87]
  PIN line[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 274.720 600.000 275.320 ;
    END
  END line[88]
  PIN line[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 277.440 600.000 278.040 ;
    END
  END line[89]
  PIN line[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 24.480 600.000 25.080 ;
    END
  END line[8]
  PIN line[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 280.840 600.000 281.440 ;
    END
  END line[90]
  PIN line[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 284.240 600.000 284.840 ;
    END
  END line[91]
  PIN line[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 286.960 600.000 287.560 ;
    END
  END line[92]
  PIN line[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 290.360 600.000 290.960 ;
    END
  END line[93]
  PIN line[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 293.080 600.000 293.680 ;
    END
  END line[94]
  PIN line[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 296.480 600.000 297.080 ;
    END
  END line[95]
  PIN line[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 299.880 600.000 300.480 ;
    END
  END line[96]
  PIN line[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 302.600 600.000 303.200 ;
    END
  END line[97]
  PIN line[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 306.000 600.000 306.600 ;
    END
  END line[98]
  PIN line[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 308.720 600.000 309.320 ;
    END
  END line[99]
  PIN line[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 27.880 600.000 28.480 ;
    END
  END line[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.440 4.000 6.040 ;
    END
  END rst_n
  PIN wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.200 4.000 10.800 ;
    END
  END wr
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 9.240 483.440 387.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 9.240 329.840 387.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 9.240 176.240 387.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 9.240 22.640 387.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 9.240 560.240 387.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 9.240 406.640 387.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 9.240 253.040 387.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 9.240 99.440 387.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 9.395 595.095 387.645 ;
      LAYER met1 ;
        RECT 5.520 9.240 595.170 388.200 ;
      LAYER met2 ;
        RECT 6.990 0.115 595.610 396.925 ;
      LAYER met3 ;
        RECT 4.000 396.760 595.600 396.905 ;
        RECT 4.400 396.040 595.600 396.760 ;
        RECT 4.400 395.360 596.000 396.040 ;
        RECT 4.000 394.040 596.000 395.360 ;
        RECT 4.000 392.640 595.600 394.040 ;
        RECT 4.000 392.000 596.000 392.640 ;
        RECT 4.400 391.320 596.000 392.000 ;
        RECT 4.400 390.600 595.600 391.320 ;
        RECT 4.000 389.920 595.600 390.600 ;
        RECT 4.000 387.920 596.000 389.920 ;
        RECT 4.000 387.240 595.600 387.920 ;
        RECT 4.400 386.520 595.600 387.240 ;
        RECT 4.400 385.840 596.000 386.520 ;
        RECT 4.000 385.200 596.000 385.840 ;
        RECT 4.000 383.800 595.600 385.200 ;
        RECT 4.000 382.480 596.000 383.800 ;
        RECT 4.400 381.800 596.000 382.480 ;
        RECT 4.400 381.080 595.600 381.800 ;
        RECT 4.000 380.400 595.600 381.080 ;
        RECT 4.000 378.400 596.000 380.400 ;
        RECT 4.000 377.720 595.600 378.400 ;
        RECT 4.400 377.000 595.600 377.720 ;
        RECT 4.400 376.320 596.000 377.000 ;
        RECT 4.000 375.680 596.000 376.320 ;
        RECT 4.000 374.280 595.600 375.680 ;
        RECT 4.000 372.960 596.000 374.280 ;
        RECT 4.400 372.280 596.000 372.960 ;
        RECT 4.400 371.560 595.600 372.280 ;
        RECT 4.000 370.880 595.600 371.560 ;
        RECT 4.000 369.560 596.000 370.880 ;
        RECT 4.000 368.200 595.600 369.560 ;
        RECT 4.400 368.160 595.600 368.200 ;
        RECT 4.400 366.800 596.000 368.160 ;
        RECT 4.000 366.160 596.000 366.800 ;
        RECT 4.000 364.760 595.600 366.160 ;
        RECT 4.000 363.440 596.000 364.760 ;
        RECT 4.400 362.760 596.000 363.440 ;
        RECT 4.400 362.040 595.600 362.760 ;
        RECT 4.000 361.360 595.600 362.040 ;
        RECT 4.000 360.040 596.000 361.360 ;
        RECT 4.000 358.680 595.600 360.040 ;
        RECT 4.400 358.640 595.600 358.680 ;
        RECT 4.400 357.280 596.000 358.640 ;
        RECT 4.000 356.640 596.000 357.280 ;
        RECT 4.000 355.240 595.600 356.640 ;
        RECT 4.000 353.920 596.000 355.240 ;
        RECT 4.400 352.520 595.600 353.920 ;
        RECT 4.000 350.520 596.000 352.520 ;
        RECT 4.000 349.160 595.600 350.520 ;
        RECT 4.400 349.120 595.600 349.160 ;
        RECT 4.400 347.760 596.000 349.120 ;
        RECT 4.000 347.120 596.000 347.760 ;
        RECT 4.000 345.720 595.600 347.120 ;
        RECT 4.000 344.400 596.000 345.720 ;
        RECT 4.400 343.000 595.600 344.400 ;
        RECT 4.000 341.000 596.000 343.000 ;
        RECT 4.000 339.640 595.600 341.000 ;
        RECT 4.400 339.600 595.600 339.640 ;
        RECT 4.400 338.280 596.000 339.600 ;
        RECT 4.400 338.240 595.600 338.280 ;
        RECT 4.000 336.880 595.600 338.240 ;
        RECT 4.000 334.880 596.000 336.880 ;
        RECT 4.400 333.480 595.600 334.880 ;
        RECT 4.000 331.480 596.000 333.480 ;
        RECT 4.000 330.120 595.600 331.480 ;
        RECT 4.400 330.080 595.600 330.120 ;
        RECT 4.400 328.760 596.000 330.080 ;
        RECT 4.400 328.720 595.600 328.760 ;
        RECT 4.000 327.360 595.600 328.720 ;
        RECT 4.000 325.360 596.000 327.360 ;
        RECT 4.400 323.960 595.600 325.360 ;
        RECT 4.000 322.640 596.000 323.960 ;
        RECT 4.000 321.240 595.600 322.640 ;
        RECT 4.000 320.600 596.000 321.240 ;
        RECT 4.400 319.240 596.000 320.600 ;
        RECT 4.400 319.200 595.600 319.240 ;
        RECT 4.000 317.840 595.600 319.200 ;
        RECT 4.000 315.840 596.000 317.840 ;
        RECT 4.400 314.440 595.600 315.840 ;
        RECT 4.000 313.120 596.000 314.440 ;
        RECT 4.000 311.720 595.600 313.120 ;
        RECT 4.000 311.080 596.000 311.720 ;
        RECT 4.400 309.720 596.000 311.080 ;
        RECT 4.400 309.680 595.600 309.720 ;
        RECT 4.000 308.320 595.600 309.680 ;
        RECT 4.000 307.000 596.000 308.320 ;
        RECT 4.000 306.320 595.600 307.000 ;
        RECT 4.400 305.600 595.600 306.320 ;
        RECT 4.400 304.920 596.000 305.600 ;
        RECT 4.000 303.600 596.000 304.920 ;
        RECT 4.000 302.200 595.600 303.600 ;
        RECT 4.000 301.560 596.000 302.200 ;
        RECT 4.400 300.880 596.000 301.560 ;
        RECT 4.400 300.160 595.600 300.880 ;
        RECT 4.000 299.480 595.600 300.160 ;
        RECT 4.000 297.480 596.000 299.480 ;
        RECT 4.000 296.800 595.600 297.480 ;
        RECT 4.400 296.080 595.600 296.800 ;
        RECT 4.400 295.400 596.000 296.080 ;
        RECT 4.000 294.080 596.000 295.400 ;
        RECT 4.000 292.680 595.600 294.080 ;
        RECT 4.000 292.040 596.000 292.680 ;
        RECT 4.400 291.360 596.000 292.040 ;
        RECT 4.400 290.640 595.600 291.360 ;
        RECT 4.000 289.960 595.600 290.640 ;
        RECT 4.000 287.960 596.000 289.960 ;
        RECT 4.000 287.280 595.600 287.960 ;
        RECT 4.400 286.560 595.600 287.280 ;
        RECT 4.400 285.880 596.000 286.560 ;
        RECT 4.000 285.240 596.000 285.880 ;
        RECT 4.000 283.840 595.600 285.240 ;
        RECT 4.000 282.520 596.000 283.840 ;
        RECT 4.400 281.840 596.000 282.520 ;
        RECT 4.400 281.120 595.600 281.840 ;
        RECT 4.000 280.440 595.600 281.120 ;
        RECT 4.000 278.440 596.000 280.440 ;
        RECT 4.000 277.760 595.600 278.440 ;
        RECT 4.400 277.040 595.600 277.760 ;
        RECT 4.400 276.360 596.000 277.040 ;
        RECT 4.000 275.720 596.000 276.360 ;
        RECT 4.000 274.320 595.600 275.720 ;
        RECT 4.000 273.000 596.000 274.320 ;
        RECT 4.400 272.320 596.000 273.000 ;
        RECT 4.400 271.600 595.600 272.320 ;
        RECT 4.000 270.920 595.600 271.600 ;
        RECT 4.000 269.600 596.000 270.920 ;
        RECT 4.000 268.240 595.600 269.600 ;
        RECT 4.400 268.200 595.600 268.240 ;
        RECT 4.400 266.840 596.000 268.200 ;
        RECT 4.000 266.200 596.000 266.840 ;
        RECT 4.000 264.800 595.600 266.200 ;
        RECT 4.000 263.480 596.000 264.800 ;
        RECT 4.400 262.800 596.000 263.480 ;
        RECT 4.400 262.080 595.600 262.800 ;
        RECT 4.000 261.400 595.600 262.080 ;
        RECT 4.000 260.080 596.000 261.400 ;
        RECT 4.000 258.720 595.600 260.080 ;
        RECT 4.400 258.680 595.600 258.720 ;
        RECT 4.400 257.320 596.000 258.680 ;
        RECT 4.000 256.680 596.000 257.320 ;
        RECT 4.000 255.280 595.600 256.680 ;
        RECT 4.000 253.960 596.000 255.280 ;
        RECT 4.400 252.560 595.600 253.960 ;
        RECT 4.000 250.560 596.000 252.560 ;
        RECT 4.000 249.200 595.600 250.560 ;
        RECT 4.400 249.160 595.600 249.200 ;
        RECT 4.400 247.800 596.000 249.160 ;
        RECT 4.000 247.160 596.000 247.800 ;
        RECT 4.000 245.760 595.600 247.160 ;
        RECT 4.000 244.440 596.000 245.760 ;
        RECT 4.400 243.040 595.600 244.440 ;
        RECT 4.000 241.040 596.000 243.040 ;
        RECT 4.000 239.680 595.600 241.040 ;
        RECT 4.400 239.640 595.600 239.680 ;
        RECT 4.400 238.320 596.000 239.640 ;
        RECT 4.400 238.280 595.600 238.320 ;
        RECT 4.000 236.920 595.600 238.280 ;
        RECT 4.000 234.920 596.000 236.920 ;
        RECT 4.400 233.520 595.600 234.920 ;
        RECT 4.000 231.520 596.000 233.520 ;
        RECT 4.000 230.160 595.600 231.520 ;
        RECT 4.400 230.120 595.600 230.160 ;
        RECT 4.400 228.800 596.000 230.120 ;
        RECT 4.400 228.760 595.600 228.800 ;
        RECT 4.000 227.400 595.600 228.760 ;
        RECT 4.000 225.400 596.000 227.400 ;
        RECT 4.400 224.000 595.600 225.400 ;
        RECT 4.000 222.680 596.000 224.000 ;
        RECT 4.000 221.280 595.600 222.680 ;
        RECT 4.000 220.640 596.000 221.280 ;
        RECT 4.400 219.280 596.000 220.640 ;
        RECT 4.400 219.240 595.600 219.280 ;
        RECT 4.000 217.880 595.600 219.240 ;
        RECT 4.000 215.880 596.000 217.880 ;
        RECT 4.400 214.480 595.600 215.880 ;
        RECT 4.000 213.160 596.000 214.480 ;
        RECT 4.000 211.760 595.600 213.160 ;
        RECT 4.000 211.120 596.000 211.760 ;
        RECT 4.400 209.760 596.000 211.120 ;
        RECT 4.400 209.720 595.600 209.760 ;
        RECT 4.000 208.360 595.600 209.720 ;
        RECT 4.000 207.040 596.000 208.360 ;
        RECT 4.000 206.360 595.600 207.040 ;
        RECT 4.400 205.640 595.600 206.360 ;
        RECT 4.400 204.960 596.000 205.640 ;
        RECT 4.000 203.640 596.000 204.960 ;
        RECT 4.000 202.240 595.600 203.640 ;
        RECT 4.000 201.600 596.000 202.240 ;
        RECT 4.400 200.920 596.000 201.600 ;
        RECT 4.400 200.200 595.600 200.920 ;
        RECT 4.000 199.520 595.600 200.200 ;
        RECT 4.000 197.520 596.000 199.520 ;
        RECT 4.000 196.840 595.600 197.520 ;
        RECT 4.400 196.120 595.600 196.840 ;
        RECT 4.400 195.440 596.000 196.120 ;
        RECT 4.000 194.120 596.000 195.440 ;
        RECT 4.000 192.720 595.600 194.120 ;
        RECT 4.000 192.080 596.000 192.720 ;
        RECT 4.400 191.400 596.000 192.080 ;
        RECT 4.400 190.680 595.600 191.400 ;
        RECT 4.000 190.000 595.600 190.680 ;
        RECT 4.000 188.000 596.000 190.000 ;
        RECT 4.000 187.320 595.600 188.000 ;
        RECT 4.400 186.600 595.600 187.320 ;
        RECT 4.400 185.920 596.000 186.600 ;
        RECT 4.000 185.280 596.000 185.920 ;
        RECT 4.000 183.880 595.600 185.280 ;
        RECT 4.000 182.560 596.000 183.880 ;
        RECT 4.400 181.880 596.000 182.560 ;
        RECT 4.400 181.160 595.600 181.880 ;
        RECT 4.000 180.480 595.600 181.160 ;
        RECT 4.000 178.480 596.000 180.480 ;
        RECT 4.000 177.800 595.600 178.480 ;
        RECT 4.400 177.080 595.600 177.800 ;
        RECT 4.400 176.400 596.000 177.080 ;
        RECT 4.000 175.760 596.000 176.400 ;
        RECT 4.000 174.360 595.600 175.760 ;
        RECT 4.000 173.040 596.000 174.360 ;
        RECT 4.400 172.360 596.000 173.040 ;
        RECT 4.400 171.640 595.600 172.360 ;
        RECT 4.000 170.960 595.600 171.640 ;
        RECT 4.000 169.640 596.000 170.960 ;
        RECT 4.000 168.280 595.600 169.640 ;
        RECT 4.400 168.240 595.600 168.280 ;
        RECT 4.400 166.880 596.000 168.240 ;
        RECT 4.000 166.240 596.000 166.880 ;
        RECT 4.000 164.840 595.600 166.240 ;
        RECT 4.000 163.520 596.000 164.840 ;
        RECT 4.400 162.840 596.000 163.520 ;
        RECT 4.400 162.120 595.600 162.840 ;
        RECT 4.000 161.440 595.600 162.120 ;
        RECT 4.000 160.120 596.000 161.440 ;
        RECT 4.000 158.760 595.600 160.120 ;
        RECT 4.400 158.720 595.600 158.760 ;
        RECT 4.400 157.360 596.000 158.720 ;
        RECT 4.000 156.720 596.000 157.360 ;
        RECT 4.000 155.320 595.600 156.720 ;
        RECT 4.000 154.000 596.000 155.320 ;
        RECT 4.400 152.600 595.600 154.000 ;
        RECT 4.000 150.600 596.000 152.600 ;
        RECT 4.000 149.240 595.600 150.600 ;
        RECT 4.400 149.200 595.600 149.240 ;
        RECT 4.400 147.840 596.000 149.200 ;
        RECT 4.000 147.200 596.000 147.840 ;
        RECT 4.000 145.800 595.600 147.200 ;
        RECT 4.000 144.480 596.000 145.800 ;
        RECT 4.400 143.080 595.600 144.480 ;
        RECT 4.000 141.080 596.000 143.080 ;
        RECT 4.000 139.720 595.600 141.080 ;
        RECT 4.400 139.680 595.600 139.720 ;
        RECT 4.400 138.360 596.000 139.680 ;
        RECT 4.400 138.320 595.600 138.360 ;
        RECT 4.000 136.960 595.600 138.320 ;
        RECT 4.000 134.960 596.000 136.960 ;
        RECT 4.400 133.560 595.600 134.960 ;
        RECT 4.000 131.560 596.000 133.560 ;
        RECT 4.000 130.200 595.600 131.560 ;
        RECT 4.400 130.160 595.600 130.200 ;
        RECT 4.400 128.840 596.000 130.160 ;
        RECT 4.400 128.800 595.600 128.840 ;
        RECT 4.000 127.440 595.600 128.800 ;
        RECT 4.000 125.440 596.000 127.440 ;
        RECT 4.400 124.040 595.600 125.440 ;
        RECT 4.000 122.720 596.000 124.040 ;
        RECT 4.000 121.320 595.600 122.720 ;
        RECT 4.000 120.680 596.000 121.320 ;
        RECT 4.400 119.320 596.000 120.680 ;
        RECT 4.400 119.280 595.600 119.320 ;
        RECT 4.000 117.920 595.600 119.280 ;
        RECT 4.000 115.920 596.000 117.920 ;
        RECT 4.400 114.520 595.600 115.920 ;
        RECT 4.000 113.200 596.000 114.520 ;
        RECT 4.000 111.800 595.600 113.200 ;
        RECT 4.000 111.160 596.000 111.800 ;
        RECT 4.400 109.800 596.000 111.160 ;
        RECT 4.400 109.760 595.600 109.800 ;
        RECT 4.000 108.400 595.600 109.760 ;
        RECT 4.000 107.080 596.000 108.400 ;
        RECT 4.000 106.400 595.600 107.080 ;
        RECT 4.400 105.680 595.600 106.400 ;
        RECT 4.400 105.000 596.000 105.680 ;
        RECT 4.000 103.680 596.000 105.000 ;
        RECT 4.000 102.280 595.600 103.680 ;
        RECT 4.000 101.640 596.000 102.280 ;
        RECT 4.400 100.960 596.000 101.640 ;
        RECT 4.400 100.240 595.600 100.960 ;
        RECT 4.000 99.560 595.600 100.240 ;
        RECT 4.000 97.560 596.000 99.560 ;
        RECT 4.000 96.880 595.600 97.560 ;
        RECT 4.400 96.160 595.600 96.880 ;
        RECT 4.400 95.480 596.000 96.160 ;
        RECT 4.000 94.160 596.000 95.480 ;
        RECT 4.000 92.760 595.600 94.160 ;
        RECT 4.000 92.120 596.000 92.760 ;
        RECT 4.400 91.440 596.000 92.120 ;
        RECT 4.400 90.720 595.600 91.440 ;
        RECT 4.000 90.040 595.600 90.720 ;
        RECT 4.000 88.040 596.000 90.040 ;
        RECT 4.000 87.360 595.600 88.040 ;
        RECT 4.400 86.640 595.600 87.360 ;
        RECT 4.400 85.960 596.000 86.640 ;
        RECT 4.000 85.320 596.000 85.960 ;
        RECT 4.000 83.920 595.600 85.320 ;
        RECT 4.000 82.600 596.000 83.920 ;
        RECT 4.400 81.920 596.000 82.600 ;
        RECT 4.400 81.200 595.600 81.920 ;
        RECT 4.000 80.520 595.600 81.200 ;
        RECT 4.000 78.520 596.000 80.520 ;
        RECT 4.000 77.840 595.600 78.520 ;
        RECT 4.400 77.120 595.600 77.840 ;
        RECT 4.400 76.440 596.000 77.120 ;
        RECT 4.000 75.800 596.000 76.440 ;
        RECT 4.000 74.400 595.600 75.800 ;
        RECT 4.000 73.080 596.000 74.400 ;
        RECT 4.400 72.400 596.000 73.080 ;
        RECT 4.400 71.680 595.600 72.400 ;
        RECT 4.000 71.000 595.600 71.680 ;
        RECT 4.000 69.680 596.000 71.000 ;
        RECT 4.000 68.320 595.600 69.680 ;
        RECT 4.400 68.280 595.600 68.320 ;
        RECT 4.400 66.920 596.000 68.280 ;
        RECT 4.000 66.280 596.000 66.920 ;
        RECT 4.000 64.880 595.600 66.280 ;
        RECT 4.000 63.560 596.000 64.880 ;
        RECT 4.400 62.880 596.000 63.560 ;
        RECT 4.400 62.160 595.600 62.880 ;
        RECT 4.000 61.480 595.600 62.160 ;
        RECT 4.000 60.160 596.000 61.480 ;
        RECT 4.000 58.800 595.600 60.160 ;
        RECT 4.400 58.760 595.600 58.800 ;
        RECT 4.400 57.400 596.000 58.760 ;
        RECT 4.000 56.760 596.000 57.400 ;
        RECT 4.000 55.360 595.600 56.760 ;
        RECT 4.000 54.040 596.000 55.360 ;
        RECT 4.400 52.640 595.600 54.040 ;
        RECT 4.000 50.640 596.000 52.640 ;
        RECT 4.000 49.280 595.600 50.640 ;
        RECT 4.400 49.240 595.600 49.280 ;
        RECT 4.400 47.880 596.000 49.240 ;
        RECT 4.000 47.240 596.000 47.880 ;
        RECT 4.000 45.840 595.600 47.240 ;
        RECT 4.000 44.520 596.000 45.840 ;
        RECT 4.400 43.120 595.600 44.520 ;
        RECT 4.000 41.120 596.000 43.120 ;
        RECT 4.000 39.760 595.600 41.120 ;
        RECT 4.400 39.720 595.600 39.760 ;
        RECT 4.400 38.400 596.000 39.720 ;
        RECT 4.400 38.360 595.600 38.400 ;
        RECT 4.000 37.000 595.600 38.360 ;
        RECT 4.000 35.000 596.000 37.000 ;
        RECT 4.400 33.600 595.600 35.000 ;
        RECT 4.000 31.600 596.000 33.600 ;
        RECT 4.000 30.240 595.600 31.600 ;
        RECT 4.400 30.200 595.600 30.240 ;
        RECT 4.400 28.880 596.000 30.200 ;
        RECT 4.400 28.840 595.600 28.880 ;
        RECT 4.000 27.480 595.600 28.840 ;
        RECT 4.000 25.480 596.000 27.480 ;
        RECT 4.400 24.080 595.600 25.480 ;
        RECT 4.000 22.760 596.000 24.080 ;
        RECT 4.000 21.360 595.600 22.760 ;
        RECT 4.000 20.720 596.000 21.360 ;
        RECT 4.400 19.360 596.000 20.720 ;
        RECT 4.400 19.320 595.600 19.360 ;
        RECT 4.000 17.960 595.600 19.320 ;
        RECT 4.000 15.960 596.000 17.960 ;
        RECT 4.400 14.560 595.600 15.960 ;
        RECT 4.000 13.240 596.000 14.560 ;
        RECT 4.000 11.840 595.600 13.240 ;
        RECT 4.000 11.200 596.000 11.840 ;
        RECT 4.400 9.840 596.000 11.200 ;
        RECT 4.400 9.800 595.600 9.840 ;
        RECT 4.000 8.440 595.600 9.800 ;
        RECT 4.000 7.120 596.000 8.440 ;
        RECT 4.000 6.440 595.600 7.120 ;
        RECT 4.400 5.720 595.600 6.440 ;
        RECT 4.400 5.040 596.000 5.720 ;
        RECT 4.000 3.720 596.000 5.040 ;
        RECT 4.000 2.320 595.600 3.720 ;
        RECT 4.000 1.680 596.000 2.320 ;
        RECT 4.400 1.000 596.000 1.680 ;
        RECT 4.400 0.280 595.600 1.000 ;
        RECT 4.000 0.135 595.600 0.280 ;
      LAYER met4 ;
        RECT 14.095 16.455 20.640 380.585 ;
        RECT 23.040 16.455 97.440 380.585 ;
        RECT 99.840 16.455 174.240 380.585 ;
        RECT 176.640 16.455 251.040 380.585 ;
        RECT 253.440 16.455 327.840 380.585 ;
        RECT 330.240 16.455 404.640 380.585 ;
        RECT 407.040 16.455 481.440 380.585 ;
        RECT 483.840 16.455 558.240 380.585 ;
        RECT 560.640 16.455 580.225 380.585 ;
  END
END DMC_32x16HC
END LIBRARY

